module redstone (tick, inputs, outputs);
	input tick;
	input [num_inputs-1:0] inputs;
	output [num_outputs:0] outputs;

parameter num_outputs = 1, num_inputs = 1;

	wire w197;
	torch #(1'b0) c197 (.i_clk(tick), .i_in(w199), .o_out(w197));
	wire w199;
	repeater #(1, 1'b0, 0, 0) c199 (.i_clk(tick), .i_in(w285), .i_lock(), .o_out(w199));
	wire w211;
	torch #(1'b1) c211 (.i_clk(tick), .i_in(w197|w224), .o_out(w211));
	wire w224;
	repeater #(1, 1'b0, 0, 0) c224 (.i_clk(tick), .i_in(w211), .i_lock(), .o_out(w224));
	wire w239;
	torch #(1'b0) c239 (.i_clk(tick), .i_in(w211), .o_out(w239));
	wire w285;
	repeater #(1, 1'b0, 0, 0) c285 (.i_clk(tick), .i_in(w350), .i_lock(), .o_out(w285));
	wire w289;
	repeater #(1, 1'b1, 0, 0) c289 (.i_clk(tick), .i_in(w239), .i_lock(), .o_out(w289));
	wire w296;
	repeater #(1, 1'b1, 0, 0) c296 (.i_clk(tick), .i_in(w239), .i_lock(), .o_out(w296));
	wire w304;
	repeater #(1, 1'b1, 1, 0) c304 (.i_clk(tick), .i_in(w289), .i_lock(), .o_out(w304));
	wire w305;
	repeater #(1, 1'b1, 0, 1) c305 (.i_clk(tick), .i_in(w306), .i_lock(w304), .o_out(w305));
	wire w306;
	repeater #(1, 1'b0, 0, 1) c306 (.i_clk(tick), .i_in(w305), .i_lock(w307), .o_out(w306));
	wire w307;
	repeater #(1, 1'b1, 1, 0) c307 (.i_clk(tick), .i_in(w296), .i_lock(), .o_out(w307));
	wire w331;
	assign outputs[0] = (w306);
	wire w350;
	assign w350 = inputs[0];
	wire w460;
	repeater #(1, 1'b1, 0, 0) c460 (.i_clk(tick), .i_in(w305), .i_lock(), .o_out(w460));
	wire w463;
	repeater #(1, 1'b1, 0, 0) c463 (.i_clk(tick), .i_in(w305), .i_lock(), .o_out(w463));
	wire w668;
	repeater #(1, 1'b1, 1, 0) c668 (.i_clk(tick), .i_in(w289|w460), .i_lock(), .o_out(w668));
	wire w669;
	repeater #(1, 1'b1, 0, 1) c669 (.i_clk(tick), .i_in(w670), .i_lock(w668), .o_out(w669));
	wire w670;
	repeater #(1, 1'b0, 0, 1) c670 (.i_clk(tick), .i_in(w669), .i_lock(w671), .o_out(w670));
	wire w671;
	repeater #(1, 1'b1, 1, 0) c671 (.i_clk(tick), .i_in(w296|w463), .i_lock(), .o_out(w671));
	wire w695;
	assign outputs[1] = (w670);
	wire w824;
	repeater #(1, 1'b1, 0, 0) c824 (.i_clk(tick), .i_in(w669), .i_lock(), .o_out(w824));
	wire w827;
	repeater #(1, 1'b1, 0, 0) c827 (.i_clk(tick), .i_in(w669), .i_lock(), .o_out(w827));
	wire w1032;
	repeater #(1, 1'b1, 1, 0) c1032 (.i_clk(tick), .i_in(w289|w460|w824), .i_lock(), .o_out(w1032));
	wire w1033;
	repeater #(1, 1'b1, 0, 1) c1033 (.i_clk(tick), .i_in(w1034), .i_lock(w1032), .o_out(w1033));
	wire w1034;
	repeater #(1, 1'b0, 0, 1) c1034 (.i_clk(tick), .i_in(w1033), .i_lock(w1035), .o_out(w1034));
	wire w1035;
	repeater #(1, 1'b1, 1, 0) c1035 (.i_clk(tick), .i_in(w296|w463|w827), .i_lock(), .o_out(w1035));
	wire w1059;
	assign outputs[2] = (w1034);
	wire w1188;
	repeater #(1, 1'b1, 0, 0) c1188 (.i_clk(tick), .i_in(w1033), .i_lock(), .o_out(w1188));
	wire w1191;
	repeater #(1, 1'b1, 0, 0) c1191 (.i_clk(tick), .i_in(w1033), .i_lock(), .o_out(w1191));
	wire w1396;
	repeater #(1, 1'b1, 1, 0) c1396 (.i_clk(tick), .i_in(w289|w460|w824|w1188), .i_lock(), .o_out(w1396));
	wire w1397;
	repeater #(1, 1'b1, 0, 1) c1397 (.i_clk(tick), .i_in(w1398), .i_lock(w1396), .o_out(w1397));
	wire w1398;
	repeater #(1, 1'b0, 0, 1) c1398 (.i_clk(tick), .i_in(w1397), .i_lock(w1399), .o_out(w1398));
	wire w1399;
	repeater #(1, 1'b1, 1, 0) c1399 (.i_clk(tick), .i_in(w296|w463|w827|w1191), .i_lock(), .o_out(w1399));
	wire w1423;
	assign outputs[3] = (w1398);
	wire w1552;
	repeater #(1, 1'b1, 0, 0) c1552 (.i_clk(tick), .i_in(w1397), .i_lock(), .o_out(w1552));
	wire w1555;
	repeater #(1, 1'b1, 0, 0) c1555 (.i_clk(tick), .i_in(w1397), .i_lock(), .o_out(w1555));
	wire w1760;
	repeater #(1, 1'b1, 1, 0) c1760 (.i_clk(tick), .i_in(w289|w460|w824|w1188|w1552), .i_lock(), .o_out(w1760));
	wire w1761;
	repeater #(1, 1'b1, 0, 1) c1761 (.i_clk(tick), .i_in(w1762), .i_lock(w1760), .o_out(w1761));
	wire w1762;
	repeater #(1, 1'b0, 0, 1) c1762 (.i_clk(tick), .i_in(w1761), .i_lock(w1763), .o_out(w1762));
	wire w1763;
	repeater #(1, 1'b1, 1, 0) c1763 (.i_clk(tick), .i_in(w296|w463|w827|w1191|w1555), .i_lock(), .o_out(w1763));
	wire w1787;
	assign outputs[4] = (w1762);
	wire w1916;
	repeater #(1, 1'b1, 0, 0) c1916 (.i_clk(tick), .i_in(w1761), .i_lock(), .o_out(w1916));
	wire w1919;
	repeater #(1, 1'b1, 0, 0) c1919 (.i_clk(tick), .i_in(w1761), .i_lock(), .o_out(w1919));
	wire w2124;
	repeater #(1, 1'b1, 1, 0) c2124 (.i_clk(tick), .i_in(w289|w460|w824|w1188|w1552|w1916), .i_lock(), .o_out(w2124));
	wire w2125;
	repeater #(1, 1'b1, 0, 1) c2125 (.i_clk(tick), .i_in(w2126), .i_lock(w2124), .o_out(w2125));
	wire w2126;
	repeater #(1, 1'b0, 0, 1) c2126 (.i_clk(tick), .i_in(w2125), .i_lock(w2127), .o_out(w2126));
	wire w2127;
	repeater #(1, 1'b1, 1, 0) c2127 (.i_clk(tick), .i_in(w296|w463|w827|w1191|w1555|w1919), .i_lock(), .o_out(w2127));
	wire w2151;
	assign outputs[5] = (w2126);
	wire w2280;
	repeater #(1, 1'b1, 0, 0) c2280 (.i_clk(tick), .i_in(w2125), .i_lock(), .o_out(w2280));
	wire w2283;
	repeater #(1, 1'b1, 0, 0) c2283 (.i_clk(tick), .i_in(w2125), .i_lock(), .o_out(w2283));
	wire w2488;
	repeater #(1, 1'b1, 1, 0) c2488 (.i_clk(tick), .i_in(w289|w460|w824|w1188|w1552|w1916|w2280), .i_lock(), .o_out(w2488));
	wire w2489;
	repeater #(1, 1'b1, 0, 1) c2489 (.i_clk(tick), .i_in(w2490), .i_lock(w2488), .o_out(w2489));
	wire w2490;
	repeater #(1, 1'b0, 0, 1) c2490 (.i_clk(tick), .i_in(w2489), .i_lock(w2491), .o_out(w2490));
	wire w2491;
	repeater #(1, 1'b1, 1, 0) c2491 (.i_clk(tick), .i_in(w296|w463|w827|w1191|w1555|w1919|w2283), .i_lock(), .o_out(w2491));
	wire w2515;
	assign outputs[6] = (w2490);
	wire w2644;
	repeater #(1, 1'b1, 0, 0) c2644 (.i_clk(tick), .i_in(w2489), .i_lock(), .o_out(w2644));
	wire w2647;
	repeater #(1, 1'b1, 0, 0) c2647 (.i_clk(tick), .i_in(w2489), .i_lock(), .o_out(w2647));
	wire w2775;
	torch #(1'b0) c2775 (.i_clk(tick), .i_in(w2814), .o_out(w2775));
	wire w2776;
	repeater #(2, 1'b1, 0, 0) c2776 (.i_clk(tick), .i_in(w2775), .i_lock(), .o_out(w2776));
	wire w2789;
	repeater #(1, 1'b0, 0, 0) c2789 (.i_clk(tick), .i_in(w2814), .i_lock(), .o_out(w2789));
	wire w2814;
	torch #(1'b1) c2814 (.i_clk(tick), .i_in(w2853), .o_out(w2814));
	wire w2852;
	repeater #(1, 1'b1, 1, 0) c2852 (.i_clk(tick), .i_in(w289|w460|w824|w1188|w1552|w1916|w2280|w2644), .i_lock(), .o_out(w2852));
	wire w2853;
	repeater #(1, 1'b1, 0, 1) c2853 (.i_clk(tick), .i_in(w2854), .i_lock(w2852), .o_out(w2853));
	wire w2854;
	repeater #(1, 1'b0, 0, 1) c2854 (.i_clk(tick), .i_in(w2853), .i_lock(w2855), .o_out(w2854));
	wire w2855;
	repeater #(1, 1'b1, 1, 0) c2855 (.i_clk(tick), .i_in(w296|w463|w827|w1191|w1555|w1919|w2283|w2647), .i_lock(), .o_out(w2855));
	wire w2879;
	assign outputs[7] = (w2854);
	wire w3201;
	repeater #(1, 1'b1, 0, 0) c3201 (.i_clk(tick), .i_in(w2776|w2789), .i_lock(), .o_out(w3201));
	wire w3208;
	repeater #(1, 1'b1, 0, 0) c3208 (.i_clk(tick), .i_in(w2776|w2789), .i_lock(), .o_out(w3208));
	wire w3216;
	repeater #(1, 1'b1, 1, 0) c3216 (.i_clk(tick), .i_in(w3201), .i_lock(), .o_out(w3216));
	wire w3217;
	repeater #(1, 1'b0, 0, 1) c3217 (.i_clk(tick), .i_in(w3218), .i_lock(w3216), .o_out(w3217));
	wire w3218;
	repeater #(1, 1'b1, 0, 1) c3218 (.i_clk(tick), .i_in(w3217), .i_lock(w3219), .o_out(w3218));
	wire w3219;
	repeater #(1, 1'b1, 1, 0) c3219 (.i_clk(tick), .i_in(w3208), .i_lock(), .o_out(w3219));
	wire w3243;
	assign outputs[8] = (w3218);
	wire w3372;
	repeater #(1, 1'b0, 0, 0) c3372 (.i_clk(tick), .i_in(w3217), .i_lock(), .o_out(w3372));
	wire w3375;
	repeater #(1, 1'b0, 0, 0) c3375 (.i_clk(tick), .i_in(w3217), .i_lock(), .o_out(w3375));
	wire w3580;
	repeater #(1, 1'b1, 1, 0) c3580 (.i_clk(tick), .i_in(w3201|w3372), .i_lock(), .o_out(w3580));
	wire w3581;
	repeater #(1, 1'b1, 0, 1) c3581 (.i_clk(tick), .i_in(w3582), .i_lock(w3580), .o_out(w3581));
	wire w3582;
	repeater #(1, 1'b0, 0, 1) c3582 (.i_clk(tick), .i_in(w3581), .i_lock(w3583), .o_out(w3582));
	wire w3583;
	repeater #(1, 1'b1, 1, 0) c3583 (.i_clk(tick), .i_in(w3208|w3375), .i_lock(), .o_out(w3583));
	wire w3607;
	assign outputs[9] = (w3582);
	wire w3736;
	repeater #(1, 1'b1, 0, 0) c3736 (.i_clk(tick), .i_in(w3581), .i_lock(), .o_out(w3736));
	wire w3739;
	repeater #(1, 1'b1, 0, 0) c3739 (.i_clk(tick), .i_in(w3581), .i_lock(), .o_out(w3739));
	wire w3944;
	repeater #(1, 1'b1, 1, 0) c3944 (.i_clk(tick), .i_in(w3201|w3372|w3736), .i_lock(), .o_out(w3944));
	wire w3945;
	repeater #(1, 1'b1, 0, 1) c3945 (.i_clk(tick), .i_in(w3946), .i_lock(w3944), .o_out(w3945));
	wire w3946;
	repeater #(1, 1'b0, 0, 1) c3946 (.i_clk(tick), .i_in(w3945), .i_lock(w3947), .o_out(w3946));
	wire w3947;
	repeater #(1, 1'b1, 1, 0) c3947 (.i_clk(tick), .i_in(w3208|w3375|w3739), .i_lock(), .o_out(w3947));
	wire w3971;
	assign outputs[10] = (w3946);
	wire w4100;
	repeater #(1, 1'b1, 0, 0) c4100 (.i_clk(tick), .i_in(w3945), .i_lock(), .o_out(w4100));
	wire w4103;
	repeater #(1, 1'b1, 0, 0) c4103 (.i_clk(tick), .i_in(w3945), .i_lock(), .o_out(w4103));
	wire w4308;
	repeater #(1, 1'b1, 1, 0) c4308 (.i_clk(tick), .i_in(w3201|w3372|w3736|w4100), .i_lock(), .o_out(w4308));
	wire w4309;
	repeater #(1, 1'b1, 0, 1) c4309 (.i_clk(tick), .i_in(w4310), .i_lock(w4308), .o_out(w4309));
	wire w4310;
	repeater #(1, 1'b0, 0, 1) c4310 (.i_clk(tick), .i_in(w4309), .i_lock(w4311), .o_out(w4310));
	wire w4311;
	repeater #(1, 1'b1, 1, 0) c4311 (.i_clk(tick), .i_in(w3208|w3375|w3739|w4103), .i_lock(), .o_out(w4311));
	wire w4335;
	assign outputs[11] = (w4310);
	wire w4464;
	repeater #(1, 1'b1, 0, 0) c4464 (.i_clk(tick), .i_in(w4309), .i_lock(), .o_out(w4464));
	wire w4467;
	repeater #(1, 1'b1, 0, 0) c4467 (.i_clk(tick), .i_in(w4309), .i_lock(), .o_out(w4467));
	wire w4672;
	repeater #(1, 1'b1, 1, 0) c4672 (.i_clk(tick), .i_in(w3201|w3372|w3736|w4100|w4464), .i_lock(), .o_out(w4672));
	wire w4673;
	repeater #(1, 1'b1, 0, 1) c4673 (.i_clk(tick), .i_in(w4674), .i_lock(w4672), .o_out(w4673));
	wire w4674;
	repeater #(1, 1'b0, 0, 1) c4674 (.i_clk(tick), .i_in(w4673), .i_lock(w4675), .o_out(w4674));
	wire w4675;
	repeater #(1, 1'b1, 1, 0) c4675 (.i_clk(tick), .i_in(w3208|w3375|w3739|w4103|w4467), .i_lock(), .o_out(w4675));
	wire w4699;
	assign outputs[12] = (w4674);
	wire w4828;
	repeater #(1, 1'b1, 0, 0) c4828 (.i_clk(tick), .i_in(w4673), .i_lock(), .o_out(w4828));
	wire w4831;
	repeater #(1, 1'b1, 0, 0) c4831 (.i_clk(tick), .i_in(w4673), .i_lock(), .o_out(w4831));
	wire w5036;
	repeater #(1, 1'b1, 1, 0) c5036 (.i_clk(tick), .i_in(w3201|w3372|w3736|w4100|w4464|w4828), .i_lock(), .o_out(w5036));
	wire w5037;
	repeater #(1, 1'b1, 0, 1) c5037 (.i_clk(tick), .i_in(w5038), .i_lock(w5036), .o_out(w5037));
	wire w5038;
	repeater #(1, 1'b0, 0, 1) c5038 (.i_clk(tick), .i_in(w5037), .i_lock(w5039), .o_out(w5038));
	wire w5039;
	repeater #(1, 1'b1, 1, 0) c5039 (.i_clk(tick), .i_in(w3208|w3375|w3739|w4103|w4467|w4831), .i_lock(), .o_out(w5039));
	wire w5063;
	assign outputs[13] = (w5038);
	wire w5192;
	repeater #(1, 1'b1, 0, 0) c5192 (.i_clk(tick), .i_in(w5037), .i_lock(), .o_out(w5192));
	wire w5195;
	repeater #(1, 1'b1, 0, 0) c5195 (.i_clk(tick), .i_in(w5037), .i_lock(), .o_out(w5195));
	wire w5400;
	repeater #(1, 1'b1, 1, 0) c5400 (.i_clk(tick), .i_in(w3201|w3372|w3736|w4100|w4464|w4828|w5192), .i_lock(), .o_out(w5400));
	wire w5401;
	repeater #(1, 1'b1, 0, 1) c5401 (.i_clk(tick), .i_in(w5402), .i_lock(w5400), .o_out(w5401));
	wire w5402;
	repeater #(1, 1'b0, 0, 1) c5402 (.i_clk(tick), .i_in(w5401), .i_lock(w5403), .o_out(w5402));
	wire w5403;
	repeater #(1, 1'b1, 1, 0) c5403 (.i_clk(tick), .i_in(w3208|w3375|w3739|w4103|w4467|w4831|w5195), .i_lock(), .o_out(w5403));
	wire w5427;
	assign outputs[14] = (w5402);
	wire w5556;
	repeater #(1, 1'b1, 0, 0) c5556 (.i_clk(tick), .i_in(w5401), .i_lock(), .o_out(w5556));
	wire w5559;
	repeater #(1, 1'b1, 0, 0) c5559 (.i_clk(tick), .i_in(w5401), .i_lock(), .o_out(w5559));
	wire w5687;
	torch #(1'b0) c5687 (.i_clk(tick), .i_in(w5726), .o_out(w5687));
	wire w5688;
	repeater #(2, 1'b1, 0, 0) c5688 (.i_clk(tick), .i_in(w5687), .i_lock(), .o_out(w5688));
	wire w5701;
	repeater #(1, 1'b0, 0, 0) c5701 (.i_clk(tick), .i_in(w5726), .i_lock(), .o_out(w5701));
	wire w5726;
	torch #(1'b1) c5726 (.i_clk(tick), .i_in(w5765), .o_out(w5726));
	wire w5764;
	repeater #(1, 1'b1, 1, 0) c5764 (.i_clk(tick), .i_in(w3201|w3372|w3736|w4100|w4464|w4828|w5192|w5556), .i_lock(), .o_out(w5764));
	wire w5765;
	repeater #(1, 1'b1, 0, 1) c5765 (.i_clk(tick), .i_in(w5766), .i_lock(w5764), .o_out(w5765));
	wire w5766;
	repeater #(1, 1'b0, 0, 1) c5766 (.i_clk(tick), .i_in(w5765), .i_lock(w5767), .o_out(w5766));
	wire w5767;
	repeater #(1, 1'b1, 1, 0) c5767 (.i_clk(tick), .i_in(w3208|w3375|w3739|w4103|w4467|w4831|w5195|w5559), .i_lock(), .o_out(w5767));
	wire w5791;
	assign outputs[15] = (w5766);
	wire w6113;
	repeater #(1, 1'b1, 0, 0) c6113 (.i_clk(tick), .i_in(w5688|w5701), .i_lock(), .o_out(w6113));
	wire w6120;
	repeater #(1, 1'b1, 0, 0) c6120 (.i_clk(tick), .i_in(w5688|w5701), .i_lock(), .o_out(w6120));
	wire w6128;
	repeater #(1, 1'b1, 1, 0) c6128 (.i_clk(tick), .i_in(w6113), .i_lock(), .o_out(w6128));
	wire w6129;
	repeater #(1, 1'b0, 0, 1) c6129 (.i_clk(tick), .i_in(w6130), .i_lock(w6128), .o_out(w6129));
	wire w6130;
	repeater #(1, 1'b1, 0, 1) c6130 (.i_clk(tick), .i_in(w6129), .i_lock(w6131), .o_out(w6130));
	wire w6131;
	repeater #(1, 1'b1, 1, 0) c6131 (.i_clk(tick), .i_in(w6120), .i_lock(), .o_out(w6131));
	wire w6155;
	assign outputs[16] = (w6130);
	wire w6284;
	repeater #(1, 1'b0, 0, 0) c6284 (.i_clk(tick), .i_in(w6129), .i_lock(), .o_out(w6284));
	wire w6287;
	repeater #(1, 1'b0, 0, 0) c6287 (.i_clk(tick), .i_in(w6129), .i_lock(), .o_out(w6287));
	wire w6492;
	repeater #(1, 1'b1, 1, 0) c6492 (.i_clk(tick), .i_in(w6113|w6284), .i_lock(), .o_out(w6492));
	wire w6493;
	repeater #(1, 1'b1, 0, 1) c6493 (.i_clk(tick), .i_in(w6494), .i_lock(w6492), .o_out(w6493));
	wire w6494;
	repeater #(1, 1'b0, 0, 1) c6494 (.i_clk(tick), .i_in(w6493), .i_lock(w6495), .o_out(w6494));
	wire w6495;
	repeater #(1, 1'b1, 1, 0) c6495 (.i_clk(tick), .i_in(w6120|w6287), .i_lock(), .o_out(w6495));
	wire w6519;
	assign outputs[17] = (w6494);
	wire w6648;
	repeater #(1, 1'b1, 0, 0) c6648 (.i_clk(tick), .i_in(w6493), .i_lock(), .o_out(w6648));
	wire w6651;
	repeater #(1, 1'b1, 0, 0) c6651 (.i_clk(tick), .i_in(w6493), .i_lock(), .o_out(w6651));
	wire w6856;
	repeater #(1, 1'b1, 1, 0) c6856 (.i_clk(tick), .i_in(w6113|w6284|w6648), .i_lock(), .o_out(w6856));
	wire w6857;
	repeater #(1, 1'b1, 0, 1) c6857 (.i_clk(tick), .i_in(w6858), .i_lock(w6856), .o_out(w6857));
	wire w6858;
	repeater #(1, 1'b0, 0, 1) c6858 (.i_clk(tick), .i_in(w6857), .i_lock(w6859), .o_out(w6858));
	wire w6859;
	repeater #(1, 1'b1, 1, 0) c6859 (.i_clk(tick), .i_in(w6120|w6287|w6651), .i_lock(), .o_out(w6859));
	wire w6883;
	assign outputs[18] = (w6858);
	wire w7012;
	repeater #(1, 1'b1, 0, 0) c7012 (.i_clk(tick), .i_in(w6857), .i_lock(), .o_out(w7012));
	wire w7015;
	repeater #(1, 1'b1, 0, 0) c7015 (.i_clk(tick), .i_in(w6857), .i_lock(), .o_out(w7015));
	wire w7220;
	repeater #(1, 1'b1, 1, 0) c7220 (.i_clk(tick), .i_in(w6113|w6284|w6648|w7012), .i_lock(), .o_out(w7220));
	wire w7221;
	repeater #(1, 1'b1, 0, 1) c7221 (.i_clk(tick), .i_in(w7222), .i_lock(w7220), .o_out(w7221));
	wire w7222;
	repeater #(1, 1'b0, 0, 1) c7222 (.i_clk(tick), .i_in(w7221), .i_lock(w7223), .o_out(w7222));
	wire w7223;
	repeater #(1, 1'b1, 1, 0) c7223 (.i_clk(tick), .i_in(w6120|w6287|w6651|w7015), .i_lock(), .o_out(w7223));
	wire w7247;
	assign outputs[19] = (w7222);
	wire w7376;
	repeater #(1, 1'b1, 0, 0) c7376 (.i_clk(tick), .i_in(w7221), .i_lock(), .o_out(w7376));
	wire w7379;
	repeater #(1, 1'b1, 0, 0) c7379 (.i_clk(tick), .i_in(w7221), .i_lock(), .o_out(w7379));
	wire w7584;
	repeater #(1, 1'b1, 1, 0) c7584 (.i_clk(tick), .i_in(w6113|w6284|w6648|w7012|w7376), .i_lock(), .o_out(w7584));
	wire w7585;
	repeater #(1, 1'b1, 0, 1) c7585 (.i_clk(tick), .i_in(w7586), .i_lock(w7584), .o_out(w7585));
	wire w7586;
	repeater #(1, 1'b0, 0, 1) c7586 (.i_clk(tick), .i_in(w7585), .i_lock(w7587), .o_out(w7586));
	wire w7587;
	repeater #(1, 1'b1, 1, 0) c7587 (.i_clk(tick), .i_in(w6120|w6287|w6651|w7015|w7379), .i_lock(), .o_out(w7587));
	wire w7611;
	assign outputs[20] = (w7586);
	wire w7740;
	repeater #(1, 1'b1, 0, 0) c7740 (.i_clk(tick), .i_in(w7585), .i_lock(), .o_out(w7740));
	wire w7743;
	repeater #(1, 1'b1, 0, 0) c7743 (.i_clk(tick), .i_in(w7585), .i_lock(), .o_out(w7743));
	wire w7948;
	repeater #(1, 1'b1, 1, 0) c7948 (.i_clk(tick), .i_in(w6113|w6284|w6648|w7012|w7376|w7740), .i_lock(), .o_out(w7948));
	wire w7949;
	repeater #(1, 1'b1, 0, 1) c7949 (.i_clk(tick), .i_in(w7950), .i_lock(w7948), .o_out(w7949));
	wire w7950;
	repeater #(1, 1'b0, 0, 1) c7950 (.i_clk(tick), .i_in(w7949), .i_lock(w7951), .o_out(w7950));
	wire w7951;
	repeater #(1, 1'b1, 1, 0) c7951 (.i_clk(tick), .i_in(w6120|w6287|w6651|w7015|w7379|w7743), .i_lock(), .o_out(w7951));
	wire w7975;
	assign outputs[21] = (w7950);
	wire w8104;
	repeater #(1, 1'b1, 0, 0) c8104 (.i_clk(tick), .i_in(w7949), .i_lock(), .o_out(w8104));
	wire w8107;
	repeater #(1, 1'b1, 0, 0) c8107 (.i_clk(tick), .i_in(w7949), .i_lock(), .o_out(w8107));
	wire w8312;
	repeater #(1, 1'b1, 1, 0) c8312 (.i_clk(tick), .i_in(w6113|w6284|w6648|w7012|w7376|w7740|w8104), .i_lock(), .o_out(w8312));
	wire w8313;
	repeater #(1, 1'b1, 0, 1) c8313 (.i_clk(tick), .i_in(w8314), .i_lock(w8312), .o_out(w8313));
	wire w8314;
	repeater #(1, 1'b0, 0, 1) c8314 (.i_clk(tick), .i_in(w8313), .i_lock(w8315), .o_out(w8314));
	wire w8315;
	repeater #(1, 1'b1, 1, 0) c8315 (.i_clk(tick), .i_in(w6120|w6287|w6651|w7015|w7379|w7743|w8107), .i_lock(), .o_out(w8315));
	wire w8339;
	assign outputs[22] = (w8314);
	wire w8468;
	repeater #(1, 1'b1, 0, 0) c8468 (.i_clk(tick), .i_in(w8313), .i_lock(), .o_out(w8468));
	wire w8471;
	repeater #(1, 1'b0, 0, 0) c8471 (.i_clk(tick), .i_in(w8313), .i_lock(), .o_out(w8471));
	wire w8599;
	torch #(1'b0) c8599 (.i_clk(tick), .i_in(w8638), .o_out(w8599));
	wire w8600;
	repeater #(2, 1'b1, 0, 0) c8600 (.i_clk(tick), .i_in(w8599), .i_lock(), .o_out(w8600));
	wire w8613;
	repeater #(1, 1'b0, 0, 0) c8613 (.i_clk(tick), .i_in(w8638), .i_lock(), .o_out(w8613));
	wire w8638;
	torch #(1'b1) c8638 (.i_clk(tick), .i_in(w8677), .o_out(w8638));
	wire w8676;
	repeater #(1, 1'b1, 1, 0) c8676 (.i_clk(tick), .i_in(w6113|w6284|w6648|w7012|w7376|w7740|w8104|w8468), .i_lock(), .o_out(w8676));
	wire w8677;
	repeater #(1, 1'b1, 0, 1) c8677 (.i_clk(tick), .i_in(w8678), .i_lock(w8676), .o_out(w8677));
	wire w8678;
	repeater #(1, 1'b0, 0, 1) c8678 (.i_clk(tick), .i_in(w8677), .i_lock(w8679), .o_out(w8678));
	wire w8679;
	repeater #(1, 1'b1, 1, 0) c8679 (.i_clk(tick), .i_in(w6120|w6287|w6651|w7015|w7379|w7743|w8107|w8471), .i_lock(), .o_out(w8679));
	wire w8703;
	assign outputs[23] = (w8678);
	wire w9025;
	repeater #(1, 1'b1, 0, 0) c9025 (.i_clk(tick), .i_in(w8600|w8613), .i_lock(), .o_out(w9025));
	wire w9032;
	repeater #(1, 1'b1, 0, 0) c9032 (.i_clk(tick), .i_in(w8600|w8613), .i_lock(), .o_out(w9032));
	wire w9040;
	repeater #(1, 1'b1, 1, 0) c9040 (.i_clk(tick), .i_in(w9025), .i_lock(), .o_out(w9040));
	wire w9041;
	repeater #(1, 1'b0, 0, 1) c9041 (.i_clk(tick), .i_in(w9042), .i_lock(w9040), .o_out(w9041));
	wire w9042;
	repeater #(1, 1'b1, 0, 1) c9042 (.i_clk(tick), .i_in(w9041), .i_lock(w9043), .o_out(w9042));
	wire w9043;
	repeater #(1, 1'b1, 1, 0) c9043 (.i_clk(tick), .i_in(w9032), .i_lock(), .o_out(w9043));
	wire w9067;
	assign outputs[24] = (w9042);
	wire w9196;
	repeater #(1, 1'b0, 0, 0) c9196 (.i_clk(tick), .i_in(w9041), .i_lock(), .o_out(w9196));
	wire w9199;
	repeater #(1, 1'b0, 0, 0) c9199 (.i_clk(tick), .i_in(w9041), .i_lock(), .o_out(w9199));
	wire w9404;
	repeater #(1, 1'b1, 1, 0) c9404 (.i_clk(tick), .i_in(w9025|w9196), .i_lock(), .o_out(w9404));
	wire w9405;
	repeater #(1, 1'b1, 0, 1) c9405 (.i_clk(tick), .i_in(w9406), .i_lock(w9404), .o_out(w9405));
	wire w9406;
	repeater #(1, 1'b0, 0, 1) c9406 (.i_clk(tick), .i_in(w9405), .i_lock(w9407), .o_out(w9406));
	wire w9407;
	repeater #(1, 1'b1, 1, 0) c9407 (.i_clk(tick), .i_in(w9032|w9199), .i_lock(), .o_out(w9407));
	wire w9431;
	assign outputs[25] = (w9406);
	wire w9560;
	repeater #(1, 1'b1, 0, 0) c9560 (.i_clk(tick), .i_in(w9405), .i_lock(), .o_out(w9560));
	wire w9563;
	repeater #(1, 1'b1, 0, 0) c9563 (.i_clk(tick), .i_in(w9405), .i_lock(), .o_out(w9563));
	wire w9768;
	repeater #(1, 1'b1, 1, 0) c9768 (.i_clk(tick), .i_in(w9025|w9196|w9560), .i_lock(), .o_out(w9768));
	wire w9769;
	repeater #(1, 1'b1, 0, 1) c9769 (.i_clk(tick), .i_in(w9770), .i_lock(w9768), .o_out(w9769));
	wire w9770;
	repeater #(1, 1'b0, 0, 1) c9770 (.i_clk(tick), .i_in(w9769), .i_lock(w9771), .o_out(w9770));
	wire w9771;
	repeater #(1, 1'b1, 1, 0) c9771 (.i_clk(tick), .i_in(w9032|w9199|w9563), .i_lock(), .o_out(w9771));
	wire w9795;
	assign outputs[26] = (w9770);
	wire w9924;
	repeater #(1, 1'b1, 0, 0) c9924 (.i_clk(tick), .i_in(w9769), .i_lock(), .o_out(w9924));
	wire w9927;
	repeater #(1, 1'b1, 0, 0) c9927 (.i_clk(tick), .i_in(w9769), .i_lock(), .o_out(w9927));
	wire w10132;
	repeater #(1, 1'b1, 1, 0) c10132 (.i_clk(tick), .i_in(w9025|w9196|w9560|w9924), .i_lock(), .o_out(w10132));
	wire w10133;
	repeater #(1, 1'b1, 0, 1) c10133 (.i_clk(tick), .i_in(w10134), .i_lock(w10132), .o_out(w10133));
	wire w10134;
	repeater #(1, 1'b0, 0, 1) c10134 (.i_clk(tick), .i_in(w10133), .i_lock(w10135), .o_out(w10134));
	wire w10135;
	repeater #(1, 1'b1, 1, 0) c10135 (.i_clk(tick), .i_in(w9032|w9199|w9563|w9927), .i_lock(), .o_out(w10135));
	wire w10159;
	assign outputs[27] = (w10134);
	wire w10288;
	repeater #(1, 1'b1, 0, 0) c10288 (.i_clk(tick), .i_in(w10133), .i_lock(), .o_out(w10288));
	wire w10291;
	repeater #(1, 1'b1, 0, 0) c10291 (.i_clk(tick), .i_in(w10133), .i_lock(), .o_out(w10291));
	wire w10496;
	repeater #(1, 1'b1, 1, 0) c10496 (.i_clk(tick), .i_in(w9025|w9196|w9560|w9924|w10288), .i_lock(), .o_out(w10496));
	wire w10497;
	repeater #(1, 1'b1, 0, 1) c10497 (.i_clk(tick), .i_in(w10498), .i_lock(w10496), .o_out(w10497));
	wire w10498;
	repeater #(1, 1'b0, 0, 1) c10498 (.i_clk(tick), .i_in(w10497), .i_lock(w10499), .o_out(w10498));
	wire w10499;
	repeater #(1, 1'b1, 1, 0) c10499 (.i_clk(tick), .i_in(w9032|w9199|w9563|w9927|w10291), .i_lock(), .o_out(w10499));
	wire w10523;
	assign outputs[28] = (w10498);
	wire w10652;
	repeater #(1, 1'b1, 0, 0) c10652 (.i_clk(tick), .i_in(w10497), .i_lock(), .o_out(w10652));
	wire w10655;
	repeater #(1, 1'b1, 0, 0) c10655 (.i_clk(tick), .i_in(w10497), .i_lock(), .o_out(w10655));
	wire w10860;
	repeater #(1, 1'b1, 1, 0) c10860 (.i_clk(tick), .i_in(w9025|w9196|w9560|w9924|w10288|w10652), .i_lock(), .o_out(w10860));
	wire w10861;
	repeater #(1, 1'b1, 0, 1) c10861 (.i_clk(tick), .i_in(w10862), .i_lock(w10860), .o_out(w10861));
	wire w10862;
	repeater #(1, 1'b0, 0, 1) c10862 (.i_clk(tick), .i_in(w10861), .i_lock(w10863), .o_out(w10862));
	wire w10863;
	repeater #(1, 1'b1, 1, 0) c10863 (.i_clk(tick), .i_in(w9032|w9199|w9563|w9927|w10291|w10655), .i_lock(), .o_out(w10863));
	wire w10887;
	assign outputs[29] = (w10862);
	wire w11016;
	repeater #(1, 1'b1, 0, 0) c11016 (.i_clk(tick), .i_in(w10861), .i_lock(), .o_out(w11016));
	wire w11019;
	repeater #(1, 1'b1, 0, 0) c11019 (.i_clk(tick), .i_in(w10861), .i_lock(), .o_out(w11019));
	wire w11224;
	repeater #(1, 1'b1, 1, 0) c11224 (.i_clk(tick), .i_in(w9025|w9196|w9560|w9924|w10288|w10652|w11016), .i_lock(), .o_out(w11224));
	wire w11225;
	repeater #(1, 1'b1, 0, 1) c11225 (.i_clk(tick), .i_in(w11226), .i_lock(w11224), .o_out(w11225));
	wire w11226;
	repeater #(1, 1'b0, 0, 1) c11226 (.i_clk(tick), .i_in(w11225), .i_lock(w11227), .o_out(w11226));
	wire w11227;
	repeater #(1, 1'b1, 1, 0) c11227 (.i_clk(tick), .i_in(w9032|w9199|w9563|w9927|w10291|w10655|w11019), .i_lock(), .o_out(w11227));
	wire w11251;
	assign outputs[30] = (w11226);
	wire w11380;
	repeater #(1, 1'b1, 0, 0) c11380 (.i_clk(tick), .i_in(w11225), .i_lock(), .o_out(w11380));
	wire w11383;
	repeater #(1, 1'b1, 0, 0) c11383 (.i_clk(tick), .i_in(w11225), .i_lock(), .o_out(w11383));
	wire w11588;
	repeater #(1, 1'b1, 1, 0) c11588 (.i_clk(tick), .i_in(w9025|w9196|w9560|w9924|w10288|w10652|w11016|w11380), .i_lock(), .o_out(w11588));
	wire w11589;
	repeater #(1, 1'b1, 0, 1) c11589 (.i_clk(tick), .i_in(w11590), .i_lock(w11588), .o_out(w11589));
	wire w11590;
	repeater #(1, 1'b0, 0, 1) c11590 (.i_clk(tick), .i_in(w11589), .i_lock(w11591), .o_out(w11590));
	wire w11591;
	repeater #(1, 1'b1, 1, 0) c11591 (.i_clk(tick), .i_in(w9032|w9199|w9563|w9927|w10291|w10655|w11019|w11383), .i_lock(), .o_out(w11591));
	wire w11615;
	assign outputs[31] = (w11590);
endmodule