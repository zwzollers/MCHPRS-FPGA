module redstone (tick, inputs, outputs);
	input tick;
	input [9:0] inputs;
	output [9:0] outputs;

	wire w60037;
	repeater #(1, 1'b0, 0, 0) c60037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60037));
	wire w64037;
	repeater #(1, 1'b0, 0, 0) c64037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64037));
	wire w68037;
	repeater #(1, 1'b0, 0, 0) c68037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68037));
	wire w72037;
	repeater #(1, 1'b0, 0, 0) c72037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72037));
	wire w76037;
	repeater #(1, 1'b0, 0, 0) c76037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76037));
	wire w80037;
	repeater #(1, 1'b0, 0, 0) c80037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80037));
	wire w84037;
	repeater #(1, 1'b0, 0, 0) c84037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84037));
	wire w60055;
	repeater #(1, 1'b0, 0, 0) c60055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60055));
	wire w64055;
	repeater #(1, 1'b0, 0, 0) c64055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64055));
	wire w68055;
	repeater #(1, 1'b0, 0, 0) c68055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68055));
	wire w72055;
	repeater #(1, 1'b0, 0, 0) c72055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72055));
	wire w76055;
	repeater #(1, 1'b0, 0, 0) c76055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76055));
	wire w80055;
	repeater #(1, 1'b0, 0, 0) c80055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80055));
	wire w84055;
	repeater #(1, 1'b0, 0, 0) c84055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84055));
	wire w70138;
	repeater #(1, 1'b0, 0, 0) c70138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70138));
	wire w54072;
	repeater #(1, 1'b0, 0, 0) c54072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54072));
	wire w42169;
	torch #(1'b0) c42169 (.i_clk(tick), .i_in(), .o_out(w42169));
	wire w46169;
	torch #(1'b0) c46169 (.i_clk(tick), .i_in(), .o_out(w46169));
	wire w50169;
	torch #(1'b0) c50169 (.i_clk(tick), .i_in(), .o_out(w50169));
	wire w54169;
	torch #(1'b0) c54169 (.i_clk(tick), .i_in(), .o_out(w54169));
	wire w58169;
	torch #(1'b0) c58169 (.i_clk(tick), .i_in(), .o_out(w58169));
	wire w62169;
	torch #(1'b0) c62169 (.i_clk(tick), .i_in(), .o_out(w62169));
	wire w66169;
	torch #(1'b0) c66169 (.i_clk(tick), .i_in(), .o_out(w66169));
	wire w29041;
	torch #(1'b0) c29041 (.i_clk(tick), .i_in(), .o_out(w29041));
	wire w33041;
	torch #(1'b0) c33041 (.i_clk(tick), .i_in(), .o_out(w33041));
	wire w37041;
	torch #(1'b0) c37041 (.i_clk(tick), .i_in(), .o_out(w37041));
	wire w41041;
	torch #(1'b0) c41041 (.i_clk(tick), .i_in(), .o_out(w41041));
	wire w45041;
	torch #(1'b0) c45041 (.i_clk(tick), .i_in(), .o_out(w45041));
	wire w49041;
	torch #(1'b0) c49041 (.i_clk(tick), .i_in(), .o_out(w49041));
	wire w53041;
	torch #(1'b0) c53041 (.i_clk(tick), .i_in(), .o_out(w53041));
	wire w57047;
	torch #(1'b1) c57047 (.i_clk(tick), .i_in(), .o_out(w57047));
	wire w58048;
	repeater #(1, 1'b0, 0, 0) c58048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58048));
	wire w60048;
	repeater #(1, 1'b1, 0, 0) c60048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60048));
	wire w62048;
	torch #(1'b1) c62048 (.i_clk(tick), .i_in(), .o_out(w62048));
	wire w28049;
	repeater #(1, 1'b0, 0, 0) c28049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28049));
	wire w32049;
	repeater #(1, 1'b0, 0, 0) c32049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32049));
	wire w36049;
	repeater #(1, 1'b0, 0, 0) c36049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36049));
	wire w40049;
	repeater #(1, 1'b0, 0, 0) c40049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40049));
	wire w44049;
	repeater #(1, 1'b0, 0, 0) c44049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44049));
	wire w48049;
	repeater #(1, 1'b0, 0, 0) c48049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48049));
	wire w52049;
	repeater #(1, 1'b0, 0, 0) c52049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52049));
	wire w56058;
	repeater #(1, 1'b1, 0, 0) c56058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56058));
	wire w28060;
	repeater #(1, 1'b0, 0, 0) c28060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28060));
	wire w32060;
	repeater #(1, 1'b0, 0, 0) c32060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32060));
	wire w36060;
	repeater #(1, 1'b0, 0, 0) c36060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36060));
	wire w40060;
	repeater #(1, 1'b0, 0, 0) c40060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40060));
	wire w44060;
	repeater #(1, 1'b0, 0, 0) c44060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44060));
	wire w48060;
	repeater #(1, 1'b0, 0, 0) c48060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48060));
	wire w52060;
	repeater #(1, 1'b0, 0, 0) c52060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52060));
	wire w57060;
	torch #(1'b1) c57060 (.i_clk(tick), .i_in(), .o_out(w57060));
	wire w29061;
	torch #(1'b0) c29061 (.i_clk(tick), .i_in(), .o_out(w29061));
	wire w33061;
	torch #(1'b0) c33061 (.i_clk(tick), .i_in(), .o_out(w33061));
	wire w37061;
	torch #(1'b0) c37061 (.i_clk(tick), .i_in(), .o_out(w37061));
	wire w41061;
	torch #(1'b0) c41061 (.i_clk(tick), .i_in(), .o_out(w41061));
	wire w45061;
	torch #(1'b0) c45061 (.i_clk(tick), .i_in(), .o_out(w45061));
	wire w49061;
	torch #(1'b0) c49061 (.i_clk(tick), .i_in(), .o_out(w49061));
	wire w53061;
	torch #(1'b0) c53061 (.i_clk(tick), .i_in(), .o_out(w53061));
	wire w58061;
	repeater #(1, 1'b0, 0, 0) c58061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58061));
	wire w62061;
	repeater #(1, 1'b1, 0, 0) c62061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62061));
	wire w56074;
	repeater #(1, 1'b1, 0, 0) c56074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56074));
	wire w28076;
	repeater #(1, 1'b0, 0, 0) c28076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28076));
	wire w32076;
	repeater #(1, 1'b0, 0, 0) c32076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32076));
	wire w36076;
	repeater #(1, 1'b0, 0, 0) c36076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36076));
	wire w40076;
	repeater #(1, 1'b0, 0, 0) c40076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40076));
	wire w44076;
	repeater #(1, 1'b0, 0, 0) c44076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44076));
	wire w48076;
	repeater #(1, 1'b0, 0, 0) c48076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48076));
	wire w52076;
	repeater #(1, 1'b0, 0, 0) c52076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52076));
	wire w57076;
	torch #(1'b0) c57076 (.i_clk(tick), .i_in(), .o_out(w57076));
	wire w29077;
	torch #(1'b0) c29077 (.i_clk(tick), .i_in(), .o_out(w29077));
	wire w33077;
	torch #(1'b0) c33077 (.i_clk(tick), .i_in(), .o_out(w33077));
	wire w37077;
	torch #(1'b0) c37077 (.i_clk(tick), .i_in(), .o_out(w37077));
	wire w41077;
	torch #(1'b0) c41077 (.i_clk(tick), .i_in(), .o_out(w41077));
	wire w45077;
	torch #(1'b0) c45077 (.i_clk(tick), .i_in(), .o_out(w45077));
	wire w49077;
	torch #(1'b0) c49077 (.i_clk(tick), .i_in(), .o_out(w49077));
	wire w53077;
	torch #(1'b0) c53077 (.i_clk(tick), .i_in(), .o_out(w53077));
	wire w58077;
	repeater #(1, 1'b0, 0, 0) c58077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58077));
	wire w56090;
	repeater #(1, 1'b0, 0, 0) c56090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56090));
	wire w28092;
	repeater #(1, 1'b0, 0, 0) c28092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28092));
	wire w32092;
	repeater #(1, 1'b0, 0, 0) c32092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32092));
	wire w36092;
	repeater #(1, 1'b0, 0, 0) c36092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36092));
	wire w40092;
	repeater #(1, 1'b0, 0, 0) c40092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40092));
	wire w44092;
	repeater #(1, 1'b0, 0, 0) c44092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44092));
	wire w48092;
	repeater #(1, 1'b0, 0, 0) c48092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48092));
	wire w52092;
	repeater #(1, 1'b0, 0, 0) c52092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52092));
	wire w57092;
	torch #(1'b1) c57092 (.i_clk(tick), .i_in(), .o_out(w57092));
	wire w73092;
	assign w73092 = inputs[0];
	wire w29093;
	torch #(1'b0) c29093 (.i_clk(tick), .i_in(), .o_out(w29093));
	wire w33093;
	torch #(1'b0) c33093 (.i_clk(tick), .i_in(), .o_out(w33093));
	wire w37093;
	torch #(1'b0) c37093 (.i_clk(tick), .i_in(), .o_out(w37093));
	wire w41093;
	torch #(1'b0) c41093 (.i_clk(tick), .i_in(), .o_out(w41093));
	wire w45093;
	torch #(1'b0) c45093 (.i_clk(tick), .i_in(), .o_out(w45093));
	wire w49093;
	torch #(1'b0) c49093 (.i_clk(tick), .i_in(), .o_out(w49093));
	wire w53093;
	torch #(1'b0) c53093 (.i_clk(tick), .i_in(), .o_out(w53093));
	wire w60093;
	repeater #(1, 1'b1, 0, 0) c60093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60093));
	wire w62093;
	repeater #(1, 1'b1, 0, 0) c62093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62093));
	wire w560106;
	repeater #(1, 1'b0, 0, 0) c560106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560106));
	wire w280108;
	repeater #(1, 1'b0, 0, 0) c280108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280108));
	wire w320108;
	repeater #(1, 1'b0, 0, 0) c320108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320108));
	wire w360108;
	repeater #(1, 1'b0, 0, 0) c360108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360108));
	wire w400108;
	repeater #(1, 1'b0, 0, 0) c400108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400108));
	wire w440108;
	repeater #(1, 1'b0, 0, 0) c440108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440108));
	wire w480108;
	repeater #(1, 1'b0, 0, 0) c480108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480108));
	wire w520108;
	repeater #(1, 1'b0, 0, 0) c520108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520108));
	wire w570108;
	torch #(1'b1) c570108 (.i_clk(tick), .i_in(), .o_out(w570108));
	wire w290109;
	torch #(1'b0) c290109 (.i_clk(tick), .i_in(), .o_out(w290109));
	wire w330109;
	torch #(1'b0) c330109 (.i_clk(tick), .i_in(), .o_out(w330109));
	wire w370109;
	torch #(1'b0) c370109 (.i_clk(tick), .i_in(), .o_out(w370109));
	wire w410109;
	torch #(1'b0) c410109 (.i_clk(tick), .i_in(), .o_out(w410109));
	wire w450109;
	torch #(1'b0) c450109 (.i_clk(tick), .i_in(), .o_out(w450109));
	wire w490109;
	torch #(1'b0) c490109 (.i_clk(tick), .i_in(), .o_out(w490109));
	wire w530109;
	torch #(1'b0) c530109 (.i_clk(tick), .i_in(), .o_out(w530109));
	wire w600109;
	repeater #(1, 1'b1, 0, 0) c600109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600109));
	wire w270112;
	repeater #(1, 1'b1, 0, 0) c270112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w270112));
	wire w280112;
	repeater #(1, 1'b0, 0, 0) c280112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280112));
	wire w310112;
	repeater #(1, 1'b1, 0, 0) c310112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310112));
	wire w320112;
	repeater #(1, 1'b0, 0, 0) c320112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320112));
	wire w350112;
	repeater #(1, 1'b1, 0, 0) c350112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w350112));
	wire w360112;
	repeater #(1, 1'b0, 0, 0) c360112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360112));
	wire w390112;
	repeater #(1, 1'b1, 0, 0) c390112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390112));
	wire w400112;
	repeater #(1, 1'b0, 0, 0) c400112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400112));
	wire w430112;
	repeater #(1, 1'b1, 0, 0) c430112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w430112));
	wire w440112;
	repeater #(1, 1'b0, 0, 0) c440112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440112));
	wire w470112;
	repeater #(1, 1'b1, 0, 0) c470112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470112));
	wire w480112;
	repeater #(1, 1'b0, 0, 0) c480112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480112));
	wire w510112;
	repeater #(1, 1'b1, 0, 0) c510112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510112));
	wire w520112;
	repeater #(1, 1'b0, 0, 0) c520112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520112));
	wire w560121;
	repeater #(4, 1'b0, 0, 0) c560121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560121));
	wire w280124;
	repeater #(1, 1'b0, 0, 0) c280124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280124));
	wire w320124;
	repeater #(1, 1'b0, 0, 0) c320124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320124));
	wire w360124;
	repeater #(1, 1'b0, 0, 0) c360124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360124));
	wire w400124;
	repeater #(1, 1'b0, 0, 0) c400124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400124));
	wire w440124;
	repeater #(1, 1'b0, 0, 0) c440124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440124));
	wire w480124;
	repeater #(1, 1'b0, 0, 0) c480124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480124));
	wire w520124;
	repeater #(1, 1'b0, 0, 0) c520124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520124));
	wire w270135;
	repeater #(1, 1'b1, 0, 0) c270135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w270135));
	wire w280135;
	repeater #(1, 1'b0, 0, 0) c280135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280135));
	wire w310135;
	repeater #(1, 1'b1, 0, 0) c310135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310135));
	wire w320135;
	repeater #(1, 1'b0, 0, 0) c320135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320135));
	wire w350135;
	repeater #(1, 1'b1, 0, 0) c350135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w350135));
	wire w360135;
	repeater #(1, 1'b0, 0, 0) c360135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360135));
	wire w390135;
	repeater #(1, 1'b1, 0, 0) c390135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390135));
	wire w400135;
	repeater #(1, 1'b0, 0, 0) c400135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400135));
	wire w430135;
	repeater #(1, 1'b1, 0, 0) c430135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w430135));
	wire w440135;
	repeater #(1, 1'b0, 0, 0) c440135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440135));
	wire w470135;
	repeater #(1, 1'b1, 0, 0) c470135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470135));
	wire w480135;
	repeater #(1, 1'b0, 0, 0) c480135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480135));
	wire w510135;
	repeater #(1, 1'b1, 0, 0) c510135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510135));
	wire w520135;
	repeater #(1, 1'b0, 0, 0) c520135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520135));
	wire w56149;
	torch #(1'b1) c56149 (.i_clk(tick), .i_in(), .o_out(w56149));
	wire w55158;
	torch #(1'b1) c55158 (.i_clk(tick), .i_in(), .o_out(w55158));
	wire w59160;
	torch #(1'b1) c59160 (.i_clk(tick), .i_in(), .o_out(w59160));
	wire w55174;
	torch #(1'b1) c55174 (.i_clk(tick), .i_in(), .o_out(w55174));
	wire w59176;
	torch #(1'b1) c59176 (.i_clk(tick), .i_in(), .o_out(w59176));
	wire w61176;
	torch #(1'b1) c61176 (.i_clk(tick), .i_in(), .o_out(w61176));
	wire w55190;
	torch #(1'b0) c55190 (.i_clk(tick), .i_in(), .o_out(w55190));
	wire w59192;
	torch #(1'b0) c59192 (.i_clk(tick), .i_in(), .o_out(w59192));
	wire w73193;
	torch #(1'b0) c73193 (.i_clk(tick), .i_in(), .o_out(w73193));
	wire w73199;
	torch #(1'b0) c73199 (.i_clk(tick), .i_in(), .o_out(w73199));
	wire w551106;
	torch #(1'b0) c551106 (.i_clk(tick), .i_in(), .o_out(w551106));
	wire w591108;
	torch #(1'b0) c591108 (.i_clk(tick), .i_in(), .o_out(w591108));
	wire w611108;
	torch #(1'b1) c611108 (.i_clk(tick), .i_in(), .o_out(w611108));
	wire w2300;
	torch #(1'b0) c2300 (.i_clk(tick), .i_in(), .o_out(w2300));
	wire w2302;
	repeater #(4, 1'b0, 0, 0) c2302 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2302));
	wire w13085;

	wire w17085;

	wire w21085;

	wire w25085;

	wire w29085;

	wire w33085;

	wire w37085;

	wire w13086;

	wire w14086;
	repeater #(2, 1'b0, 0, 0) c14086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14086));
	wire w17086;

	wire w18086;
	repeater #(2, 1'b0, 0, 0) c18086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18086));
	wire w21086;

	wire w22086;
	repeater #(2, 1'b0, 0, 0) c22086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22086));
	wire w25086;

	wire w26086;
	repeater #(2, 1'b0, 0, 0) c26086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26086));
	wire w29086;

	wire w30086;
	repeater #(2, 1'b0, 0, 0) c30086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30086));
	wire w33086;

	wire w34086;
	repeater #(2, 1'b0, 0, 0) c34086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34086));
	wire w37086;

	wire w38086;
	repeater #(2, 1'b0, 0, 0) c38086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38086));
	wire w41086;
	repeater #(2, 1'b0, 0, 0) c41086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41086));
	wire w13087;
	repeater #(1, 1'b0, 0, 0) c13087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13087));
	wire w17087;
	repeater #(1, 1'b0, 0, 0) c17087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17087));
	wire w21087;
	repeater #(1, 1'b0, 0, 0) c21087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21087));
	wire w25087;
	repeater #(1, 1'b0, 0, 0) c25087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25087));
	wire w29087;
	repeater #(1, 1'b0, 0, 0) c29087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29087));
	wire w33087;
	repeater #(1, 1'b0, 0, 0) c33087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33087));
	wire w37087;
	repeater #(1, 1'b0, 0, 0) c37087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37087));
	wire w40089;
	repeater #(2, 1'b0, 0, 0) c40089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40089));
	wire w40091;
	torch #(1'b1) c40091 (.i_clk(tick), .i_in(), .o_out(w40091));
	wire w130101;
	repeater #(1, 1'b1, 0, 0) c130101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130101));
	wire w170101;
	repeater #(1, 1'b1, 0, 0) c170101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170101));
	wire w210101;
	repeater #(1, 1'b1, 0, 0) c210101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210101));
	wire w250101;
	repeater #(1, 1'b1, 0, 0) c250101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250101));
	wire w290101;
	repeater #(2, 1'b1, 0, 0) c290101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290101));
	wire w330101;
	repeater #(2, 1'b1, 0, 0) c330101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330101));
	wire w370101;
	repeater #(2, 1'b1, 0, 0) c370101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370101));
	wire w400101;
	repeater #(1, 1'b1, 0, 0) c400101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400101));
	wire w420101;
	repeater #(1, 1'b0, 0, 0) c420101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420101));
	wire w440101;
	repeater #(1, 1'b1, 0, 0) c440101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440101));
	wire w460101;
	repeater #(1, 1'b1, 0, 0) c460101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460101));
	wire w130102;
	repeater #(1, 1'b0, 0, 0) c130102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130102));
	wire w140102;
	repeater #(1, 1'b0, 0, 0) c140102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140102));
	wire w170102;
	repeater #(1, 1'b0, 0, 0) c170102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170102));
	wire w180102;
	repeater #(1, 1'b0, 0, 0) c180102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180102));
	wire w210102;
	repeater #(1, 1'b0, 0, 0) c210102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210102));
	wire w220102;
	repeater #(1, 1'b0, 0, 0) c220102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220102));
	wire w250102;
	repeater #(1, 1'b0, 0, 0) c250102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250102));
	wire w260102;
	repeater #(1, 1'b0, 0, 0) c260102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260102));
	wire w290102;
	repeater #(1, 1'b0, 0, 0) c290102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290102));
	wire w300102;
	repeater #(1, 1'b0, 0, 0) c300102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300102));
	wire w330102;
	repeater #(1, 1'b0, 0, 0) c330102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330102));
	wire w340102;
	repeater #(1, 1'b0, 0, 0) c340102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340102));
	wire w370102;
	repeater #(1, 1'b0, 0, 0) c370102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370102));
	wire w130103;

	wire w170103;

	wire w210103;

	wire w250103;

	wire w290103;

	wire w330103;

	wire w370103;

	wire w230106;
	torch #(1'b1) c230106 (.i_clk(tick), .i_in(), .o_out(w230106));
	wire w360108;
	repeater #(1, 1'b1, 0, 0) c360108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360108));
	wire w810110;
	repeater #(1, 1'b0, 0, 0) c810110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w810110));
	wire w1150110;
	repeater #(1, 1'b0, 0, 0) c1150110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1150110));
	wire w130117;
	repeater #(1, 1'b1, 0, 0) c130117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130117));
	wire w170117;
	repeater #(1, 1'b1, 0, 0) c170117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170117));
	wire w210117;
	repeater #(1, 1'b1, 0, 0) c210117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210117));
	wire w250117;
	repeater #(1, 1'b1, 0, 0) c250117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250117));
	wire w290117;
	repeater #(2, 1'b1, 0, 0) c290117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290117));
	wire w330117;
	repeater #(2, 1'b1, 0, 0) c330117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330117));
	wire w370117;
	repeater #(2, 1'b1, 0, 0) c370117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370117));
	wire w400117;
	repeater #(1, 1'b1, 0, 0) c400117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400117));
	wire w420117;
	repeater #(1, 1'b0, 0, 0) c420117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420117));
	wire w440117;
	repeater #(1, 1'b1, 0, 0) c440117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440117));
	wire w460117;
	repeater #(1, 1'b1, 0, 0) c460117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460117));
	wire w130118;
	repeater #(1, 1'b0, 0, 0) c130118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130118));
	wire w140118;
	repeater #(1, 1'b0, 0, 0) c140118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140118));
	wire w170118;
	repeater #(1, 1'b0, 0, 0) c170118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170118));
	wire w180118;
	repeater #(1, 1'b0, 0, 0) c180118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180118));
	wire w210118;
	repeater #(1, 1'b0, 0, 0) c210118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210118));
	wire w220118;
	repeater #(1, 1'b0, 0, 0) c220118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220118));
	wire w250118;
	repeater #(1, 1'b0, 0, 0) c250118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250118));
	wire w260118;
	repeater #(1, 1'b0, 0, 0) c260118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260118));
	wire w290118;
	repeater #(1, 1'b0, 0, 0) c290118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290118));
	wire w300118;
	repeater #(1, 1'b0, 0, 0) c300118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300118));
	wire w330118;
	repeater #(1, 1'b0, 0, 0) c330118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330118));
	wire w340118;
	repeater #(1, 1'b0, 0, 0) c340118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340118));
	wire w370118;
	repeater #(1, 1'b0, 0, 0) c370118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370118));
	wire w130119;

	wire w170119;

	wire w210119;

	wire w250119;

	wire w290119;

	wire w330119;

	wire w370119;

	wire w230122;
	torch #(1'b1) c230122 (.i_clk(tick), .i_in(), .o_out(w230122));
	wire w360124;
	repeater #(1, 1'b1, 0, 0) c360124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360124));
	wire w570126;

	wire w560127;

	wire w580127;

	wire w560129;

	wire w580129;

	wire w560131;

	wire w580131;

	wire w130133;
	repeater #(1, 1'b1, 0, 0) c130133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130133));
	wire w170133;
	repeater #(1, 1'b1, 0, 0) c170133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170133));
	wire w210133;
	repeater #(1, 1'b1, 0, 0) c210133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210133));
	wire w250133;
	repeater #(1, 1'b1, 0, 0) c250133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250133));
	wire w290133;
	repeater #(2, 1'b1, 0, 0) c290133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290133));
	wire w330133;
	repeater #(2, 1'b1, 0, 0) c330133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330133));
	wire w370133;
	repeater #(2, 1'b1, 0, 0) c370133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370133));
	wire w400133;
	repeater #(1, 1'b1, 0, 0) c400133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400133));
	wire w420133;
	repeater #(1, 1'b0, 0, 0) c420133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420133));
	wire w440133;
	repeater #(1, 1'b1, 0, 0) c440133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440133));
	wire w460133;
	repeater #(1, 1'b1, 0, 0) c460133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460133));
	wire w560133;

	wire w580133;

	wire w130134;
	repeater #(1, 1'b0, 0, 0) c130134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130134));
	wire w140134;
	repeater #(1, 1'b0, 0, 0) c140134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140134));
	wire w170134;
	repeater #(1, 1'b0, 0, 0) c170134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170134));
	wire w180134;
	repeater #(1, 1'b0, 0, 0) c180134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180134));
	wire w210134;
	repeater #(1, 1'b0, 0, 0) c210134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210134));
	wire w220134;
	repeater #(1, 1'b0, 0, 0) c220134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220134));
	wire w250134;
	repeater #(1, 1'b0, 0, 0) c250134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250134));
	wire w260134;
	repeater #(1, 1'b0, 0, 0) c260134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260134));
	wire w290134;
	repeater #(1, 1'b0, 0, 0) c290134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290134));
	wire w300134;
	repeater #(1, 1'b0, 0, 0) c300134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300134));
	wire w330134;
	repeater #(1, 1'b0, 0, 0) c330134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330134));
	wire w340134;
	repeater #(1, 1'b0, 0, 0) c340134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340134));
	wire w370134;
	repeater #(1, 1'b0, 0, 0) c370134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370134));
	wire w130135;

	wire w170135;

	wire w210135;

	wire w250135;

	wire w290135;

	wire w330135;

	wire w370135;

	wire w560135;

	wire w580135;

	wire w550137;
	repeater #(1, 1'b0, 0, 0) c550137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550137));
	wire w560137;

	wire w570137;
	repeater #(1, 1'b1, 0, 0) c570137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570137));
	wire w580137;

	wire w590137;
	repeater #(1, 1'b0, 0, 0) c590137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590137));
	wire w230138;
	torch #(1'b1) c230138 (.i_clk(tick), .i_in(), .o_out(w230138));
	wire w570138;

	wire w550139;
	repeater #(1, 1'b0, 0, 0) c550139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550139));
	wire w560139;

	wire w580139;

	wire w590139;
	repeater #(1, 1'b0, 0, 0) c590139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590139));
	wire w360140;
	repeater #(1, 1'b1, 0, 0) c360140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360140));
	wire w570140;

	wire w560141;

	wire w570141;
	repeater #(1, 1'b1, 0, 0) c570141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570141));
	wire w580141;

	wire w560143;

	wire w580143;

	wire w560145;

	wire w580145;

	wire w520146;
	repeater #(1, 1'b0, 0, 0) c520146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520146));
	wire w560147;

	wire w580147;

	wire w130149;
	repeater #(1, 1'b1, 0, 0) c130149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130149));
	wire w170149;
	repeater #(1, 1'b1, 0, 0) c170149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170149));
	wire w210149;
	repeater #(1, 1'b1, 0, 0) c210149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210149));
	wire w250149;
	repeater #(1, 1'b1, 0, 0) c250149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250149));
	wire w290149;
	repeater #(2, 1'b1, 0, 0) c290149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290149));
	wire w330149;
	repeater #(2, 1'b1, 0, 0) c330149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330149));
	wire w370149;
	repeater #(2, 1'b1, 0, 0) c370149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370149));
	wire w400149;
	repeater #(1, 1'b1, 0, 0) c400149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400149));
	wire w420149;
	repeater #(1, 1'b0, 0, 0) c420149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420149));
	wire w440149;
	repeater #(1, 1'b1, 0, 0) c440149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440149));
	wire w460149;
	repeater #(1, 1'b1, 0, 0) c460149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460149));
	wire w560149;

	wire w580149;

	wire w130150;
	repeater #(1, 1'b0, 0, 0) c130150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130150));
	wire w140150;
	repeater #(1, 1'b0, 0, 0) c140150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140150));
	wire w170150;
	repeater #(1, 1'b0, 0, 0) c170150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170150));
	wire w180150;
	repeater #(1, 1'b0, 0, 0) c180150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180150));
	wire w210150;
	repeater #(1, 1'b0, 0, 0) c210150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210150));
	wire w220150;
	repeater #(1, 1'b0, 0, 0) c220150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220150));
	wire w250150;
	repeater #(1, 1'b0, 0, 0) c250150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250150));
	wire w260150;
	repeater #(1, 1'b0, 0, 0) c260150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260150));
	wire w290150;
	repeater #(1, 1'b0, 0, 0) c290150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290150));
	wire w300150;
	repeater #(1, 1'b0, 0, 0) c300150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300150));
	wire w330150;
	repeater #(1, 1'b0, 0, 0) c330150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330150));
	wire w340150;
	repeater #(1, 1'b0, 0, 0) c340150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340150));
	wire w370150;
	repeater #(1, 1'b0, 0, 0) c370150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370150));
	wire w130151;

	wire w170151;

	wire w210151;

	wire w250151;

	wire w290151;

	wire w330151;

	wire w370151;

	wire w560151;

	wire w580151;

	wire w560153;

	wire w580153;

	wire w230154;
	torch #(1'b1) c230154 (.i_clk(tick), .i_in(), .o_out(w230154));
	wire w560155;

	wire w580155;

	wire w360156;
	repeater #(1, 1'b1, 0, 0) c360156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360156));
	wire w560157;

	wire w580157;

	wire w230159;

	wire w560159;

	wire w580159;

	wire w190160;

	wire w220160;

	wire w240160;

	wire w270160;

	wire w180161;

	wire w200161;

	wire w230161;

	wire w260161;

	wire w280161;

	wire w300161;

	wire w560161;

	wire w580161;

	wire w270162;

	wire w180163;

	wire w200163;

	wire w220163;

	wire w260163;

	wire w270163;

	wire w310163;

	wire w400163;
	repeater #(1, 1'b1, 0, 0) c400163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400163));
	wire w420163;
	repeater #(1, 1'b0, 0, 0) c420163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420163));
	wire w440163;
	repeater #(1, 1'b1, 0, 0) c440163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440163));
	wire w460163;
	repeater #(1, 1'b1, 0, 0) c460163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460163));
	wire w560163;

	wire w580163;

	wire w260164;

	wire w560165;

	wire w580165;

	wire w210166;
	repeater #(1, 1'b0, 0, 0) c210166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210166));
	wire w240166;
	repeater #(1, 1'b0, 0, 0) c240166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240166));
	wire w250166;
	repeater #(1, 1'b0, 0, 0) c250166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250166));
	wire w200167;

	wire w240167;

	wire w400167;
	repeater #(3, 1'b0, 0, 0) c400167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400167));
	wire w560167;

	wire w580167;

	wire w280169;
	torch #(1'b0) c280169 (.i_clk(tick), .i_in(), .o_out(w280169));
	wire w560169;

	wire w580169;

	wire w300170;
	torch #(1'b1) c300170 (.i_clk(tick), .i_in(), .o_out(w300170));
	wire w580171;
	repeater #(4, 1'b0, 0, 0) c580171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580171));
	wire w400173;
	repeater #(1, 1'b0, 0, 0) c400173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400173));
	wire w580173;
	repeater #(4, 1'b0, 0, 0) c580173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580173));
	wire w580175;
	repeater #(4, 1'b0, 0, 0) c580175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580175));
	wire w350177;
	assign w350177 = inputs[1];
	wire w450177;
	repeater #(1, 1'b0, 0, 0) c450177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w450177));
	wire w580177;
	repeater #(4, 1'b0, 0, 0) c580177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580177));
	wire w5610;
	repeater #(1, 1'b0, 0, 0) c5610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5610));
	wire w2311;
	repeater #(1, 1'b0, 0, 0) c2311 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2311));
	wire w5811;
	repeater #(1, 1'b0, 0, 0) c5811 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5811));
	wire w78194;

	wire w112194;

	wire w80197;

	wire w114197;

	wire w39199;
	repeater #(1, 1'b0, 0, 0) c39199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39199));
	wire w271100;
	repeater #(1, 1'b1, 0, 0) c271100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w271100));
	wire w811100;

	wire w1151100;

	wire w411101;

	wire w391103;
	torch #(1'b0) c391103 (.i_clk(tick), .i_in(), .o_out(w391103));
	wire w791103;

	wire w811103;

	wire w1131103;

	wire w1151103;

	wire w381105;
	torch #(1'b1) c381105 (.i_clk(tick), .i_in(), .o_out(w381105));
	wire w811105;

	wire w821105;

	wire w831105;

	wire w1151105;

	wire w1161105;

	wire w1171105;

	wire w381106;
	repeater #(1, 1'b0, 0, 0) c381106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w381106));
	wire w831106;

	wire w1171106;

	wire w351107;
	repeater #(1, 1'b0, 0, 0) c351107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w351107));
	wire w811108;
	repeater #(1, 1'b0, 0, 0) c811108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811108));
	wire w831108;
	torch #(1'b0) c831108 (.i_clk(tick), .i_in(), .o_out(w831108));
	wire w1151108;
	repeater #(1, 1'b0, 0, 0) c1151108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1151108));
	wire w1171108;
	torch #(1'b0) c1171108 (.i_clk(tick), .i_in(), .o_out(w1171108));
	wire w851110;
	repeater #(1, 1'b0, 0, 0) c851110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w851110));
	wire w1191110;
	repeater #(1, 1'b0, 0, 0) c1191110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1191110));
	wire w821112;
	torch #(1'b1) c821112 (.i_clk(tick), .i_in(), .o_out(w821112));
	wire w1161112;
	torch #(1'b1) c1161112 (.i_clk(tick), .i_in(), .o_out(w1161112));
	wire w391115;
	repeater #(1, 1'b0, 0, 0) c391115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w391115));
	wire w271116;
	repeater #(1, 1'b1, 0, 0) c271116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w271116));
	wire w411117;

	wire w391119;
	torch #(1'b0) c391119 (.i_clk(tick), .i_in(), .o_out(w391119));
	wire w381121;
	torch #(1'b1) c381121 (.i_clk(tick), .i_in(), .o_out(w381121));
	wire w381122;
	repeater #(1, 1'b0, 0, 0) c381122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w381122));
	wire w351123;
	repeater #(1, 1'b0, 0, 0) c351123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w351123));
	wire w391131;
	repeater #(1, 1'b0, 0, 0) c391131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w391131));
	wire w271132;
	repeater #(1, 1'b1, 0, 0) c271132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w271132));
	wire w411133;

	wire w391135;
	torch #(1'b1) c391135 (.i_clk(tick), .i_in(), .o_out(w391135));
	wire w2201;
	torch #(1'b1) c2201 (.i_clk(tick), .i_in(), .o_out(w2201));
	wire w2202;
	repeater #(1, 1'b0, 0, 0) c2202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2202));
	wire w1903;
	repeater #(1, 1'b0, 0, 0) c1903 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1903));
	wire w23011;
	repeater #(1, 1'b0, 0, 0) c23011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23011));
	wire w11012;
	repeater #(1, 1'b1, 0, 0) c11012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11012));
	wire w25013;

	wire w23015;
	torch #(1'b1) c23015 (.i_clk(tick), .i_in(), .o_out(w23015));
	wire w22017;
	torch #(1'b1) c22017 (.i_clk(tick), .i_in(), .o_out(w22017));
	wire w22018;
	repeater #(1, 1'b0, 0, 0) c22018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22018));
	wire w19019;
	repeater #(1, 1'b0, 0, 0) c19019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19019));
	wire w6030;
	repeater #(1, 1'b0, 0, 0) c6030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6030));
	wire w7030;
	repeater #(1, 1'b0, 0, 0) c7030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7030));
	wire w10030;
	repeater #(1, 1'b0, 0, 0) c10030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10030));
	wire w11030;
	repeater #(1, 1'b0, 0, 0) c11030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11030));
	wire w24030;
	torch #(1'b0) c24030 (.i_clk(tick), .i_in(), .o_out(w24030));
	wire w6031;

	wire w10031;

	wire w38032;
	torch #(1'b1) c38032 (.i_clk(tick), .i_in(), .o_out(w38032));
	wire w20033;
	repeater #(4, 1'b0, 0, 0) c20033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20033));
	wire w39034;
	repeater #(4, 1'b0, 0, 0) c39034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39034));
	wire w44034;
	repeater #(1, 1'b0, 0, 0) c44034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44034));
	wire w20035;
	repeater #(4, 1'b0, 0, 0) c20035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20035));
	wire w28035;
	torch #(1'b0) c28035 (.i_clk(tick), .i_in(), .o_out(w28035));
	wire w30035;
	torch #(1'b0) c30035 (.i_clk(tick), .i_in(), .o_out(w30035));
	wire w37035;

	wire w38035;
	repeater #(1, 1'b0, 0, 0) c38035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38035));
	wire w16036;

	wire w35036;
	repeater #(2, 1'b0, 0, 0) c35036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35036));
	wire w36036;
	repeater #(4, 1'b0, 0, 0) c36036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36036));
	wire w20037;
	repeater #(4, 1'b0, 0, 0) c20037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20037));
	wire w26037;
	torch #(1'b1) c26037 (.i_clk(tick), .i_in(), .o_out(w26037));
	wire w33037;
	repeater #(1, 1'b0, 0, 0) c33037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33037));
	wire w16038;

	wire w34038;
	repeater #(1, 1'b0, 0, 0) c34038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34038));
	wire w37038;

	wire w38038;
	repeater #(1, 1'b0, 0, 0) c38038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38038));
	wire w44038;
	repeater #(3, 1'b0, 0, 0) c44038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44038));
	wire w45038;
	torch #(1'b0) c45038 (.i_clk(tick), .i_in(), .o_out(w45038));
	wire w19039;
	repeater #(1, 1'b0, 0, 0) c19039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19039));
	wire w20039;
	repeater #(4, 1'b0, 0, 0) c20039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20039));
	wire w26039;
	torch #(1'b1) c26039 (.i_clk(tick), .i_in(), .o_out(w26039));
	wire w30039;
	torch #(1'b1) c30039 (.i_clk(tick), .i_in(), .o_out(w30039));
	wire w36039;
	repeater #(3, 1'b0, 0, 0) c36039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36039));
	wire w44039;

	wire w16040;
	repeater #(1, 1'b0, 0, 0) c16040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16040));
	wire w22041;
	torch #(1'b0) c22041 (.i_clk(tick), .i_in(), .o_out(w22041));
	wire w34041;
	repeater #(1, 1'b0, 0, 0) c34041 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34041));
	wire w37041;

	wire w38041;
	repeater #(1, 1'b0, 0, 0) c38041 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38041));
	wire w36042;
	repeater #(2, 1'b0, 0, 0) c36042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36042));
	wire w21043;
	repeater #(4, 1'b0, 0, 0) c21043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21043));
	wire w30043;
	repeater #(1, 1'b0, 0, 0) c30043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30043));
	wire w880112;
	torch #(1'b1) c880112 (.i_clk(tick), .i_in(), .o_out(w880112));
	wire w1220112;
	torch #(1'b1) c1220112 (.i_clk(tick), .i_in(), .o_out(w1220112));
	wire w870117;

	wire w1210117;

	wire w620134;

	wire w660134;

	wire w960134;

	wire w1000134;

	wire w660137;

	wire w1000137;

	wire w690139;

	wire w1030139;

	wire w260143;
	repeater #(1, 1'b1, 0, 0) c260143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260143));
	wire w690143;

	wire w1030143;

	wire w240144;
	repeater #(1, 1'b0, 0, 0) c240144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240144));
	wire w670146;

	wire w690146;

	wire w1010146;

	wire w1030146;

	wire w690148;

	wire w700148;

	wire w710148;

	wire w1030148;

	wire w1040148;

	wire w1050148;

	wire w640149;

	wire w650149;

	wire w710149;

	wire w980149;

	wire w990149;

	wire w1050149;

	wire w690151;
	repeater #(1, 1'b0, 0, 0) c690151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w690151));
	wire w710151;
	torch #(1'b0) c710151 (.i_clk(tick), .i_in(), .o_out(w710151));
	wire w1030151;
	repeater #(1, 1'b0, 0, 0) c1030151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030151));
	wire w1050151;
	torch #(1'b0) c1050151 (.i_clk(tick), .i_in(), .o_out(w1050151));
	wire w730153;
	repeater #(1, 1'b1, 0, 0) c730153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w730153));
	wire w1070153;
	repeater #(1, 1'b1, 0, 0) c1070153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070153));
	wire w700155;
	torch #(1'b1) c700155 (.i_clk(tick), .i_in(), .o_out(w700155));
	wire w1040155;
	torch #(1'b1) c1040155 (.i_clk(tick), .i_in(), .o_out(w1040155));
	wire w650158;
	repeater #(1, 1'b0, 0, 0) c650158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650158));
	wire w990158;
	repeater #(1, 1'b0, 0, 0) c990158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990158));
	wire w260159;
	repeater #(1, 1'b1, 0, 0) c260159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260159));
	wire w240160;
	repeater #(1, 1'b0, 0, 0) c240160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240160));
	wire w400168;
	repeater #(1, 1'b0, 0, 0) c400168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400168));
	wire w420168;
	repeater #(1, 1'b0, 0, 0) c420168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420168));
	wire w400172;
	repeater #(1, 1'b0, 0, 0) c400172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400172));
	wire w420172;
	repeater #(1, 1'b0, 0, 0) c420172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420172));
	wire w260175;
	repeater #(1, 1'b1, 0, 0) c260175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260175));
	wire w240176;
	repeater #(1, 1'b0, 0, 0) c240176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240176));
	wire w400176;
	repeater #(1, 1'b0, 0, 0) c400176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400176));
	wire w420176;
	repeater #(1, 1'b0, 0, 0) c420176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420176));
	wire w4011;
	repeater #(1, 1'b0, 0, 0) c4011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4011));
	wire w4211;
	repeater #(1, 1'b0, 0, 0) c4211 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4211));
	wire w4015;
	repeater #(1, 1'b0, 0, 0) c4015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4015));
	wire w4215;
	repeater #(1, 1'b0, 0, 0) c4215 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4215));
	wire w4019;
	repeater #(1, 1'b0, 0, 0) c4019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4019));
	wire w4219;
	repeater #(1, 1'b0, 0, 0) c4219 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4219));
	wire w26112;
	repeater #(1, 1'b1, 0, 0) c26112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26112));
	wire w24113;
	repeater #(1, 1'b0, 0, 0) c24113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24113));
	wire w40113;
	repeater #(1, 1'b0, 0, 0) c40113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40113));
	wire w42113;
	repeater #(1, 1'b0, 0, 0) c42113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42113));
	wire w40117;
	repeater #(1, 1'b0, 0, 0) c40117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40117));
	wire w42117;
	repeater #(1, 1'b0, 0, 0) c42117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42117));
	wire w40121;
	repeater #(1, 1'b0, 0, 0) c40121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40121));
	wire w42121;
	repeater #(1, 1'b0, 0, 0) c42121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42121));
	wire w40125;
	repeater #(1, 1'b0, 0, 0) c40125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40125));
	wire w42125;
	repeater #(1, 1'b0, 0, 0) c42125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42125));
	wire w26126;
	torch #(1'b0) c26126 (.i_clk(tick), .i_in(), .o_out(w26126));
	wire w25128;
	torch #(1'b1) c25128 (.i_clk(tick), .i_in(), .o_out(w25128));
	wire w40129;
	repeater #(1, 1'b0, 0, 0) c40129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40129));
	wire w42129;
	repeater #(1, 1'b0, 0, 0) c42129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42129));
	wire w25131;
	repeater #(1, 1'b0, 0, 0) c25131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25131));
	wire w12133;
	torch #(1'b0) c12133 (.i_clk(tick), .i_in(), .o_out(w12133));
	wire w17136;
	torch #(1'b1) c17136 (.i_clk(tick), .i_in(), .o_out(w17136));
	wire w37136;
	torch #(1'b1) c37136 (.i_clk(tick), .i_in(), .o_out(w37136));
	wire w15137;
	repeater #(2, 1'b0, 0, 0) c15137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15137));
	wire w17138;
	torch #(1'b0) c17138 (.i_clk(tick), .i_in(), .o_out(w17138));
	wire w37139;
	torch #(1'b0) c37139 (.i_clk(tick), .i_in(), .o_out(w37139));
	wire w17140;
	torch #(1'b0) c17140 (.i_clk(tick), .i_in(), .o_out(w17140));
	wire w37142;
	torch #(1'b0) c37142 (.i_clk(tick), .i_in(), .o_out(w37142));
	wire w20144;
	repeater #(1, 1'b0, 0, 0) c20144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20144));
	wire w841112;
	torch #(1'b1) c841112 (.i_clk(tick), .i_in(), .o_out(w841112));
	wire w1181112;
	torch #(1'b1) c1181112 (.i_clk(tick), .i_in(), .o_out(w1181112));
	wire w831117;

	wire w1171117;

	wire w861121;

	wire w1201121;

	wire w701134;

	wire w1041134;

	wire w4300;
	repeater #(1, 1'b1, 0, 0) c4300 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4300));
	wire w7700;
	repeater #(1, 1'b1, 0, 0) c7700 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7700));
	wire w5401;

	wire w8801;

	wire w4303;

	wire w7703;

	wire w5604;

	wire w9004;

	wire w4307;

	wire w4407;

	wire w5707;

	wire w7707;

	wire w7807;

	wire w9107;

	wire w708;
	repeater #(1, 1'b1, 0, 0) c708 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w708));
	wire w4409;

	wire w7809;

	wire w55010;

	wire w57010;

	wire w89010;

	wire w91010;

	wire w6012;
	repeater #(2, 1'b1, 0, 0) c6012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6012));
	wire w57012;

	wire w58012;

	wire w59012;

	wire w91012;

	wire w92012;

	wire w93012;

	wire w52013;

	wire w53013;

	wire w59013;

	wire w86013;

	wire w87013;

	wire w93013;

	wire w49015;
	torch #(1'b0) c49015 (.i_clk(tick), .i_in(), .o_out(w49015));
	wire w57015;
	repeater #(1, 1'b1, 0, 0) c57015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57015));
	wire w59015;
	torch #(1'b0) c59015 (.i_clk(tick), .i_in(), .o_out(w59015));
	wire w83015;
	torch #(1'b0) c83015 (.i_clk(tick), .i_in(), .o_out(w83015));
	wire w91015;
	repeater #(1, 1'b1, 0, 0) c91015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91015));
	wire w93015;
	torch #(1'b0) c93015 (.i_clk(tick), .i_in(), .o_out(w93015));
	wire w61017;
	repeater #(1, 1'b1, 0, 0) c61017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61017));
	wire w95017;
	repeater #(1, 1'b1, 0, 0) c95017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95017));
	wire w58019;
	torch #(1'b1) c58019 (.i_clk(tick), .i_in(), .o_out(w58019));
	wire w92019;
	torch #(1'b1) c92019 (.i_clk(tick), .i_in(), .o_out(w92019));
	wire w50021;
	torch #(1'b1) c50021 (.i_clk(tick), .i_in(), .o_out(w50021));
	wire w84021;
	torch #(1'b1) c84021 (.i_clk(tick), .i_in(), .o_out(w84021));
	wire w53022;
	repeater #(1, 1'b0, 0, 0) c53022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53022));
	wire w87022;
	repeater #(1, 1'b0, 0, 0) c87022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87022));
	wire w7024;
	repeater #(1, 1'b1, 0, 0) c7024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7024));
	wire w6028;
	repeater #(2, 1'b1, 0, 0) c6028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6028));
	wire w7040;
	repeater #(1, 1'b1, 0, 0) c7040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7040));
	wire w6044;
	repeater #(2, 1'b1, 0, 0) c6044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6044));
	wire w26046;
	repeater #(1, 1'b0, 0, 0) c26046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26046));
	wire w28050;
	repeater #(2, 1'b0, 0, 0) c28050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28050));
	wire w28051;

	wire w7056;
	repeater #(1, 1'b1, 0, 0) c7056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7056));
	wire w26058;
	repeater #(1, 1'b0, 0, 0) c26058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26058));
	wire w6060;
	repeater #(2, 1'b1, 0, 0) c6060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6060));
	wire w6071;
	torch #(1'b0) c6071 (.i_clk(tick), .i_in(), .o_out(w6071));
	wire w4072;
	torch #(1'b1) c4072 (.i_clk(tick), .i_in(), .o_out(w4072));
	wire w198072;
	repeater #(1, 1'b0, 0, 0) c198072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198072));
	wire w199072;
	repeater #(1, 1'b0, 0, 0) c199072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199072));
	wire w202072;
	repeater #(1, 1'b0, 0, 0) c202072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202072));
	wire w203072;
	repeater #(1, 1'b0, 0, 0) c203072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203072));
	wire w206072;
	repeater #(2, 1'b0, 0, 0) c206072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206072));
	wire w198073;

	wire w202073;

	wire w6074;
	repeater #(2, 1'b0, 0, 0) c6074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6074));
	wire w16077;
	repeater #(1, 1'b1, 0, 0) c16077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16077));
	wire w19078;
	repeater #(1, 1'b1, 0, 0) c19078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19078));
	wire w15079;
	torch #(1'b0) c15079 (.i_clk(tick), .i_in(), .o_out(w15079));
	wire w19079;
	repeater #(1, 1'b1, 0, 0) c19079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19079));
	wire w206080;
	repeater #(2, 1'b0, 0, 0) c206080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206080));
	wire w15081;
	torch #(1'b1) c15081 (.i_clk(tick), .i_in(), .o_out(w15081));
	wire w19081;
	repeater #(1, 1'b1, 0, 0) c19081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19081));
	wire w19082;
	repeater #(1, 1'b0, 0, 0) c19082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19082));
	wire w15083;
	torch #(1'b1) c15083 (.i_clk(tick), .i_in(), .o_out(w15083));
	wire w19084;
	repeater #(1, 1'b1, 0, 0) c19084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19084));
	wire w19085;
	repeater #(1, 1'b0, 0, 0) c19085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19085));
	wire w720153;
	repeater #(2, 1'b1, 0, 0) c720153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w720153));
	wire w1060153;
	repeater #(2, 1'b1, 0, 0) c1060153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060153));
	wire w640155;
	torch #(1'b0) c640155 (.i_clk(tick), .i_in(), .o_out(w640155));
	wire w740155;
	repeater #(1, 1'b1, 0, 0) c740155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w740155));
	wire w980155;
	torch #(1'b0) c980155 (.i_clk(tick), .i_in(), .o_out(w980155));
	wire w1080155;
	repeater #(1, 1'b1, 0, 0) c1080155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1080155));
	wire w740159;
	repeater #(1, 1'b1, 0, 0) c740159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w740159));
	wire w1080159;
	repeater #(1, 1'b1, 0, 0) c1080159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1080159));
	wire w630160;

	wire w970160;

	wire w740162;

	wire w1080162;

	wire w660164;

	wire w1000164;

	wire w720165;

	wire w730165;

	wire w1060165;

	wire w1070165;

	wire w660166;

	wire w700166;

	wire w1000166;

	wire w1040166;

	wire w460175;

	wire w500175;

	wire w540175;

	wire w580175;

	wire w800175;

	wire w840175;

	wire w880175;

	wire w920175;

	wire w580177;

	wire w920177;

	wire w4710;
	repeater #(1, 1'b1, 0, 0) c4710 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4710));
	wire w8110;
	repeater #(1, 1'b1, 0, 0) c8110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8110));
	wire w5811;

	wire w9211;

	wire w4713;

	wire w6113;

	wire w8113;

	wire w9513;

	wire w5814;

	wire w9214;

	wire w5515;

	wire w8915;

	wire w4717;

	wire w4817;

	wire w6117;

	wire w8117;

	wire w8217;

	wire w9517;

	wire w1018;
	repeater #(1, 1'b0, 0, 0) c1018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1018));
	wire w4819;

	wire w8219;

	wire w59110;

	wire w61110;

	wire w93110;

	wire w95110;

	wire w61112;

	wire w62112;

	wire w63112;

	wire w95112;

	wire w96112;

	wire w97112;

	wire w56113;

	wire w57113;

	wire w63113;

	wire w90113;

	wire w91113;

	wire w97113;

	wire w53115;
	torch #(1'b0) c53115 (.i_clk(tick), .i_in(), .o_out(w53115));
	wire w61115;
	repeater #(1, 1'b1, 0, 0) c61115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61115));
	wire w63115;
	torch #(1'b0) c63115 (.i_clk(tick), .i_in(), .o_out(w63115));
	wire w87115;
	torch #(1'b0) c87115 (.i_clk(tick), .i_in(), .o_out(w87115));
	wire w95115;
	repeater #(1, 1'b1, 0, 0) c95115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95115));
	wire w97115;
	torch #(1'b0) c97115 (.i_clk(tick), .i_in(), .o_out(w97115));
	wire w31117;
	assign w31117 = inputs[2];
	wire w49117;
	repeater #(1, 1'b1, 0, 0) c49117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49117));
	wire w65117;
	repeater #(1, 1'b1, 0, 0) c65117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65117));
	wire w83117;
	repeater #(1, 1'b1, 0, 0) c83117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83117));
	wire w99117;
	repeater #(1, 1'b1, 0, 0) c99117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99117));
	wire w17118;
	assign w17118 = inputs[3];
	wire w20118;
	assign w20118 = inputs[4];
	wire w62119;
	torch #(1'b1) c62119 (.i_clk(tick), .i_in(), .o_out(w62119));
	wire w96119;
	torch #(1'b1) c96119 (.i_clk(tick), .i_in(), .o_out(w96119));
	wire w54121;
	torch #(1'b1) c54121 (.i_clk(tick), .i_in(), .o_out(w54121));
	wire w88121;
	torch #(1'b1) c88121 (.i_clk(tick), .i_in(), .o_out(w88121));
	wire w57122;
	repeater #(1, 1'b0, 0, 0) c57122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57122));
	wire w91122;
	repeater #(1, 1'b0, 0, 0) c91122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91122));
	wire w51123;
	repeater #(1, 1'b0, 0, 0) c51123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51123));
	wire w85123;
	repeater #(1, 1'b0, 0, 0) c85123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85123));
	wire w10124;
	repeater #(1, 1'b0, 0, 0) c10124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10124));
	wire w51125;
	repeater #(1, 1'b0, 0, 0) c51125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51125));
	wire w85125;
	repeater #(1, 1'b0, 0, 0) c85125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85125));
	wire w10140;
	repeater #(1, 1'b0, 0, 0) c10140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10140));
	wire w10156;
	repeater #(1, 1'b0, 0, 0) c10156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10156));
	wire w23158;
	repeater #(1, 1'b0, 0, 0) c23158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23158));
	wire w4167;
	repeater #(1, 1'b0, 0, 0) c4167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4167));
	wire w5167;
	repeater #(4, 1'b0, 0, 0) c5167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5167));
	wire w4168;

	wire w4169;
	repeater #(4, 1'b0, 0, 0) c4169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4169));
	wire w10169;
	torch #(1'b1) c10169 (.i_clk(tick), .i_in(), .o_out(w10169));
	wire w21169;
	repeater #(1, 1'b0, 0, 0) c21169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21169));
	wire w9171;
	repeater #(4, 1'b1, 0, 0) c9171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9171));
	wire w9172;
	repeater #(4, 1'b1, 0, 0) c9172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9172));
	wire w9173;
	repeater #(4, 1'b1, 0, 0) c9173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9173));
	wire w23174;
	repeater #(1, 1'b0, 0, 0) c23174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23174));
	wire w12176;
	torch #(1'b0) c12176 (.i_clk(tick), .i_in(), .o_out(w12176));
	wire w6177;
	torch #(1'b0) c6177 (.i_clk(tick), .i_in(), .o_out(w6177));
	wire w205178;
	torch #(1'b1) c205178 (.i_clk(tick), .i_in(), .o_out(w205178));
	wire w0179;
	repeater #(3, 1'b0, 0, 0) c0179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0179));
	wire w205180;
	torch #(1'b1) c205180 (.i_clk(tick), .i_in(), .o_out(w205180));
	wire w0181;
	repeater #(3, 1'b1, 0, 0) c0181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0181));
	wire w205182;
	torch #(1'b1) c205182 (.i_clk(tick), .i_in(), .o_out(w205182));
	wire w0183;
	repeater #(3, 1'b1, 0, 0) c0183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0183));
	wire w52017;
	repeater #(2, 1'b1, 0, 0) c52017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52017));
	wire w86017;
	repeater #(2, 1'b1, 0, 0) c86017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86017));
	wire w44019;
	torch #(1'b0) c44019 (.i_clk(tick), .i_in(), .o_out(w44019));
	wire w54019;
	repeater #(1, 1'b1, 0, 0) c54019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54019));
	wire w78019;
	torch #(1'b0) c78019 (.i_clk(tick), .i_in(), .o_out(w78019));
	wire w88019;
	repeater #(1, 1'b1, 0, 0) c88019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88019));
	wire w54023;
	repeater #(1, 1'b1, 0, 0) c54023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54023));
	wire w88023;
	repeater #(1, 1'b1, 0, 0) c88023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88023));
	wire w43024;

	wire w77024;

	wire w54026;

	wire w88026;

	wire w43027;

	wire w77027;

	wire w46028;

	wire w80028;

	wire w52029;

	wire w53029;

	wire w86029;

	wire w87029;

	wire w46030;

	wire w80030;

	wire w30032;

	wire w34032;

	wire w38032;

	wire w42032;

	wire w46032;

	wire w50032;

	wire w54032;

	wire w64032;

	wire w68032;

	wire w72032;

	wire w76032;

	wire w80032;

	wire w84032;

	wire w88032;

	wire w30036;

	wire w34036;

	wire w38036;

	wire w42036;

	wire w46036;

	wire w50036;

	wire w54036;

	wire w64036;

	wire w68036;

	wire w72036;

	wire w76036;

	wire w80036;

	wire w84036;

	wire w88036;

	wire w28038;
	repeater #(1, 1'b1, 0, 0) c28038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28038));
	wire w32038;
	repeater #(1, 1'b1, 0, 0) c32038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32038));
	wire w36038;
	repeater #(1, 1'b1, 0, 0) c36038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36038));
	wire w40038;
	repeater #(1, 1'b0, 0, 0) c40038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40038));
	wire w62038;
	repeater #(1, 1'b1, 0, 0) c62038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62038));
	wire w66038;
	repeater #(1, 1'b1, 0, 0) c66038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66038));
	wire w70038;
	repeater #(1, 1'b0, 0, 0) c70038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70038));
	wire w74038;
	repeater #(1, 1'b1, 0, 0) c74038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74038));
	wire w46039;

	wire w50039;

	wire w54039;

	wire w80039;

	wire w84039;

	wire w88039;

	wire w46041;

	wire w80041;

	wire w35043;
	repeater #(1, 1'b1, 0, 0) c35043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35043));
	wire w69043;
	repeater #(1, 1'b0, 0, 0) c69043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69043));
	wire w30044;

	wire w46044;

	wire w64044;

	wire w80044;

	wire w38045;

	wire w72045;

	wire w33046;

	wire w35046;

	wire w41046;

	wire w49046;

	wire w67046;

	wire w69046;

	wire w75046;

	wire w83046;

	wire w46047;

	wire w80047;

	wire w205047;
	repeater #(1, 1'b0, 0, 0) c205047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205047));
	wire w206047;
	torch #(1'b0) c206047 (.i_clk(tick), .i_in(), .o_out(w206047));
	wire w43048;

	wire w44048;

	wire w77048;

	wire w78048;

	wire w206049;
	repeater #(4, 1'b0, 0, 0) c206049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206049));
	wire w33050;

	wire w35050;

	wire w36050;

	wire w49050;

	wire w67050;

	wire w69050;

	wire w70050;

	wire w83050;

	wire w30052;
	torch #(1'b1) c30052 (.i_clk(tick), .i_in(), .o_out(w30052));
	wire w31052;

	wire w36052;

	wire w64052;
	torch #(1'b1) c64052 (.i_clk(tick), .i_in(), .o_out(w64052));
	wire w65052;

	wire w70052;

	wire w31053;

	wire w33053;

	wire w47053;

	wire w49053;

	wire w65053;

	wire w67053;

	wire w81053;

	wire w83053;

	wire w33055;

	wire w34055;

	wire w35055;

	wire w49055;

	wire w50055;

	wire w51055;

	wire w67055;

	wire w68055;

	wire w69055;

	wire w83055;

	wire w84055;

	wire w85055;

	wire w35056;

	wire w44056;

	wire w45056;

	wire w51056;

	wire w69056;

	wire w78056;

	wire w79056;

	wire w85056;

	wire w33058;
	repeater #(1, 1'b0, 0, 0) c33058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33058));
	wire w35058;
	torch #(1'b0) c35058 (.i_clk(tick), .i_in(), .o_out(w35058));
	wire w41058;
	torch #(1'b1) c41058 (.i_clk(tick), .i_in(), .o_out(w41058));
	wire w49058;
	repeater #(1, 1'b1, 0, 0) c49058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49058));
	wire w51058;
	torch #(1'b0) c51058 (.i_clk(tick), .i_in(), .o_out(w51058));
	wire w67058;
	repeater #(1, 1'b0, 0, 0) c67058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67058));
	wire w69058;
	torch #(1'b0) c69058 (.i_clk(tick), .i_in(), .o_out(w69058));
	wire w75058;
	torch #(1'b1) c75058 (.i_clk(tick), .i_in(), .o_out(w75058));
	wire w83058;
	repeater #(1, 1'b1, 0, 0) c83058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83058));
	wire w85058;
	torch #(1'b0) c85058 (.i_clk(tick), .i_in(), .o_out(w85058));
	wire w2059;

	wire w37060;
	repeater #(1, 1'b1, 0, 0) c37060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37060));
	wire w53060;
	repeater #(1, 1'b0, 0, 0) c53060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53060));
	wire w71060;
	repeater #(1, 1'b1, 0, 0) c71060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71060));
	wire w87060;
	repeater #(1, 1'b0, 0, 0) c87060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87060));
	wire w34062;
	torch #(1'b1) c34062 (.i_clk(tick), .i_in(), .o_out(w34062));
	wire w50062;
	torch #(1'b1) c50062 (.i_clk(tick), .i_in(), .o_out(w50062));
	wire w68062;
	torch #(1'b1) c68062 (.i_clk(tick), .i_in(), .o_out(w68062));
	wire w84062;
	torch #(1'b1) c84062 (.i_clk(tick), .i_in(), .o_out(w84062));
	wire w206062;
	repeater #(1, 1'b0, 0, 0) c206062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206062));
	wire w42064;
	torch #(1'b1) c42064 (.i_clk(tick), .i_in(), .o_out(w42064));
	wire w76064;
	torch #(1'b1) c76064 (.i_clk(tick), .i_in(), .o_out(w76064));
	wire w33065;
	repeater #(1, 1'b0, 0, 0) c33065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33065));
	wire w45065;
	repeater #(1, 1'b0, 0, 0) c45065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45065));
	wire w67065;
	repeater #(1, 1'b0, 0, 0) c67065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67065));
	wire w79065;
	repeater #(1, 1'b0, 0, 0) c79065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79065));
	wire w39066;
	repeater #(1, 1'b0, 0, 0) c39066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39066));
	wire w73066;
	repeater #(1, 1'b0, 0, 0) c73066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73066));
	wire w39068;
	repeater #(1, 1'b0, 0, 0) c39068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39068));
	wire w73068;
	repeater #(1, 1'b0, 0, 0) c73068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73068));
	wire w172069;
	repeater #(2, 1'b0, 0, 0) c172069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172069));
	wire w176069;
	repeater #(2, 1'b0, 0, 0) c176069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176069));
	wire w180069;
	repeater #(2, 1'b0, 0, 0) c180069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180069));
	wire w184069;
	repeater #(2, 1'b0, 0, 0) c184069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184069));
	wire w188069;
	repeater #(2, 1'b0, 0, 0) c188069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188069));
	wire w192069;
	repeater #(2, 1'b0, 0, 0) c192069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192069));
	wire w196069;
	repeater #(2, 1'b0, 0, 0) c196069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196069));
	wire w172070;
	repeater #(2, 1'b0, 0, 0) c172070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172070));
	wire w176070;
	repeater #(2, 1'b0, 0, 0) c176070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176070));
	wire w180070;
	repeater #(2, 1'b0, 0, 0) c180070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180070));
	wire w184070;
	repeater #(2, 1'b0, 0, 0) c184070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184070));
	wire w188070;
	repeater #(2, 1'b0, 0, 0) c188070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188070));
	wire w192070;
	repeater #(2, 1'b0, 0, 0) c192070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192070));
	wire w196070;
	repeater #(2, 1'b0, 0, 0) c196070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196070));
	wire w206071;
	repeater #(1, 1'b0, 0, 0) c206071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206071));
	wire w206076;
	repeater #(1, 1'b0, 0, 0) c206076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206076));
	wire w172085;
	repeater #(2, 1'b0, 0, 0) c172085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172085));
	wire w176085;
	repeater #(2, 1'b0, 0, 0) c176085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176085));
	wire w180085;
	repeater #(2, 1'b0, 0, 0) c180085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180085));
	wire w184085;
	repeater #(2, 1'b0, 0, 0) c184085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184085));
	wire w188085;
	repeater #(2, 1'b0, 0, 0) c188085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188085));
	wire w192085;
	repeater #(2, 1'b0, 0, 0) c192085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192085));
	wire w196085;
	repeater #(2, 1'b0, 0, 0) c196085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196085));
	wire w175086;
	assign w175086 = inputs[5];
	wire w206087;
	repeater #(1, 1'b0, 0, 0) c206087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206087));
	wire w13095;
	repeater #(1, 1'b0, 0, 0) c13095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13095));
	wire w206097;
	repeater #(4, 1'b0, 0, 0) c206097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206097));
	wire w206098;
	repeater #(4, 1'b0, 0, 0) c206098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206098));
	wire w206099;
	repeater #(4, 1'b0, 0, 0) c206099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206099));
	wire w2060100;
	repeater #(4, 1'b0, 0, 0) c2060100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060100));
	wire w2060101;
	repeater #(4, 1'b0, 0, 0) c2060101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060101));
	wire w2060102;
	repeater #(4, 1'b0, 0, 0) c2060102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060102));
	wire w2060103;
	repeater #(4, 1'b0, 0, 0) c2060103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060103));
	wire w2060104;
	repeater #(4, 1'b0, 0, 0) c2060104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060104));
	wire w2060105;
	repeater #(4, 1'b0, 0, 0) c2060105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060105));
	wire w2060106;
	repeater #(4, 1'b0, 0, 0) c2060106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060106));
	wire w2060107;
	repeater #(4, 1'b0, 0, 0) c2060107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060107));
	wire w2060108;
	repeater #(4, 1'b0, 0, 0) c2060108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060108));
	wire w2060109;
	assign outputs[0] = ();
	wire w2060110;
	repeater #(4, 1'b0, 0, 0) c2060110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060110));
	wire w2060111;
	repeater #(4, 1'b0, 0, 0) c2060111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060111));
	wire w2060112;
	repeater #(4, 1'b0, 0, 0) c2060112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060112));
	wire w2060113;
	repeater #(4, 1'b0, 0, 0) c2060113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060113));
	wire w2060114;
	repeater #(4, 1'b0, 0, 0) c2060114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060114));
	wire w2020115;
	torch #(1'b1) c2020115 (.i_clk(tick), .i_in(), .o_out(w2020115));
	wire w2060115;
	repeater #(4, 1'b0, 0, 0) c2060115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060115));
	wire w2060116;
	repeater #(4, 1'b0, 0, 0) c2060116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060116));
	wire w2060117;
	repeater #(4, 1'b0, 0, 0) c2060117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060117));
	wire w2060118;
	repeater #(4, 1'b0, 0, 0) c2060118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060118));
	wire w2060119;
	repeater #(4, 1'b0, 0, 0) c2060119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060119));
	wire w2060120;
	repeater #(4, 1'b0, 0, 0) c2060120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060120));
	wire w1910121;
	torch #(1'b0) c1910121 (.i_clk(tick), .i_in(), .o_out(w1910121));
	wire w2060121;
	repeater #(4, 1'b0, 0, 0) c2060121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060121));
	wire w2060122;
	repeater #(4, 1'b0, 0, 0) c2060122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060122));
	wire w1910123;
	torch #(1'b1) c1910123 (.i_clk(tick), .i_in(), .o_out(w1910123));
	wire w2060123;
	repeater #(4, 1'b0, 0, 0) c2060123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060123));
	wire w1910125;
	torch #(1'b1) c1910125 (.i_clk(tick), .i_in(), .o_out(w1910125));
	wire w48117;
	repeater #(2, 1'b0, 0, 0) c48117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48117));
	wire w82117;
	repeater #(2, 1'b0, 0, 0) c82117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82117));
	wire w40119;
	torch #(1'b0) c40119 (.i_clk(tick), .i_in(), .o_out(w40119));
	wire w50119;
	repeater #(1, 1'b1, 0, 0) c50119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50119));
	wire w56119;
	torch #(1'b1) c56119 (.i_clk(tick), .i_in(), .o_out(w56119));
	wire w74119;
	torch #(1'b0) c74119 (.i_clk(tick), .i_in(), .o_out(w74119));
	wire w84119;
	repeater #(1, 1'b0, 0, 0) c84119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84119));
	wire w90119;
	torch #(1'b1) c90119 (.i_clk(tick), .i_in(), .o_out(w90119));
	wire w50123;
	repeater #(1, 1'b1, 0, 0) c50123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50123));
	wire w84123;
	repeater #(1, 1'b0, 0, 0) c84123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84123));
	wire w39124;

	wire w55124;

	wire w73124;

	wire w89124;

	wire w47125;

	wire w81125;

	wire w44126;

	wire w50126;

	wire w78126;

	wire w84126;

	wire w39127;

	wire w73127;

	wire w42128;

	wire w76128;

	wire w48129;

	wire w49129;

	wire w82129;

	wire w83129;

	wire w34130;

	wire w38130;

	wire w42130;

	wire w68130;

	wire w72130;

	wire w76130;

	wire w58133;

	wire w92133;

	wire w31134;

	wire w32134;

	wire w35134;

	wire w36134;

	wire w39134;

	wire w40134;

	wire w43134;

	wire w44134;

	wire w47134;

	wire w48134;

	wire w51134;

	wire w52134;

	wire w55134;

	wire w56134;

	wire w65134;

	wire w66134;

	wire w69134;

	wire w70134;

	wire w73134;

	wire w74134;

	wire w77134;

	wire w78134;

	wire w81134;

	wire w82134;

	wire w85134;

	wire w86134;

	wire w89134;

	wire w90134;

	wire w29135;

	wire w63135;

	wire w44138;
	repeater #(1, 1'b1, 0, 0) c44138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44138));
	wire w48138;
	repeater #(1, 1'b1, 0, 0) c48138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48138));
	wire w52138;
	repeater #(1, 1'b1, 0, 0) c52138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52138));
	wire w78138;
	repeater #(1, 1'b0, 0, 0) c78138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78138));
	wire w82138;
	repeater #(1, 1'b1, 0, 0) c82138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82138));
	wire w86138;
	repeater #(1, 1'b1, 0, 0) c86138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86138));
	wire w176138;
	repeater #(1, 1'b0, 0, 0) c176138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176138));
	wire w180138;
	repeater #(2, 1'b0, 0, 0) c180138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180138));
	wire w184138;
	repeater #(2, 1'b0, 0, 0) c184138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184138));
	wire w188138;
	repeater #(2, 1'b0, 0, 0) c188138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188138));
	wire w192138;
	repeater #(2, 1'b0, 0, 0) c192138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192138));
	wire w196138;
	repeater #(2, 1'b0, 0, 0) c196138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196138));
	wire w184139;
	repeater #(1, 1'b0, 0, 0) c184139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184139));
	wire w188139;
	repeater #(2, 1'b0, 0, 0) c188139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188139));
	wire w192139;
	repeater #(2, 1'b0, 0, 0) c192139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192139));
	wire w196139;
	repeater #(2, 1'b0, 0, 0) c196139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196139));
	wire w192140;
	repeater #(1, 1'b0, 0, 0) c192140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192140));
	wire w196140;
	repeater #(2, 1'b0, 0, 0) c196140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196140));
	wire w30141;

	wire w34141;

	wire w50141;

	wire w54141;

	wire w64141;

	wire w68141;

	wire w84141;

	wire w88141;

	wire w39143;
	repeater #(1, 1'b0, 0, 0) c39143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39143));
	wire w73143;
	repeater #(1, 1'b1, 0, 0) c73143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73143));
	wire w202143;
	repeater #(1, 1'b1, 0, 0) c202143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202143));
	wire w204143;
	repeater #(1, 1'b1, 0, 0) c204143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204143));
	wire w206143;
	repeater #(1, 1'b1, 0, 0) c206143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206143));
	wire w34144;

	wire w50144;

	wire w68144;

	wire w84144;

	wire w42145;

	wire w76145;

	wire w37146;

	wire w39146;

	wire w40146;

	wire w45146;

	wire w53146;

	wire w71146;

	wire w73146;

	wire w74146;

	wire w79146;

	wire w87146;

	wire w50147;

	wire w84147;

	wire w47148;

	wire w48148;

	wire w81148;

	wire w82148;

	wire w37150;

	wire w39150;

	wire w40150;

	wire w53150;

	wire w71150;

	wire w73150;

	wire w74150;

	wire w87150;

	wire w34152;
	torch #(1'b1) c34152 (.i_clk(tick), .i_in(), .o_out(w34152));
	wire w35152;

	wire w40152;

	wire w68152;
	torch #(1'b1) c68152 (.i_clk(tick), .i_in(), .o_out(w68152));
	wire w69152;

	wire w74152;

	wire w35153;

	wire w37153;

	wire w51153;

	wire w53153;

	wire w69153;

	wire w71153;

	wire w85153;

	wire w87153;

	wire w172154;
	repeater #(2, 1'b0, 0, 0) c172154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172154));
	wire w176154;
	repeater #(2, 1'b0, 0, 0) c176154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176154));
	wire w180154;
	repeater #(2, 1'b0, 0, 0) c180154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180154));
	wire w184154;
	repeater #(2, 1'b0, 0, 0) c184154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184154));
	wire w188154;
	repeater #(2, 1'b0, 0, 0) c188154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188154));
	wire w192154;
	repeater #(2, 1'b0, 0, 0) c192154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192154));
	wire w196154;
	repeater #(2, 1'b0, 0, 0) c196154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196154));
	wire w37155;

	wire w38155;

	wire w39155;

	wire w53155;

	wire w54155;

	wire w55155;

	wire w71155;

	wire w72155;

	wire w73155;

	wire w87155;

	wire w88155;

	wire w89155;

	wire w172155;
	repeater #(2, 1'b0, 0, 0) c172155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172155));
	wire w176155;
	repeater #(2, 1'b0, 0, 0) c176155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176155));
	wire w180155;
	repeater #(2, 1'b0, 0, 0) c180155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180155));
	wire w184155;
	repeater #(2, 1'b0, 0, 0) c184155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184155));
	wire w188155;
	repeater #(2, 1'b0, 0, 0) c188155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188155));
	wire w192155;
	repeater #(2, 1'b0, 0, 0) c192155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192155));
	wire w196155;
	repeater #(2, 1'b0, 0, 0) c196155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196155));
	wire w32156;

	wire w33156;

	wire w39156;

	wire w48156;

	wire w49156;

	wire w55156;

	wire w66156;

	wire w67156;

	wire w73156;

	wire w82156;

	wire w83156;

	wire w89156;

	wire w172156;
	repeater #(2, 1'b0, 0, 0) c172156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172156));
	wire w176156;
	repeater #(2, 1'b0, 0, 0) c176156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176156));
	wire w180156;
	repeater #(2, 1'b0, 0, 0) c180156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180156));
	wire w184156;
	repeater #(2, 1'b0, 0, 0) c184156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184156));
	wire w188156;
	repeater #(2, 1'b0, 0, 0) c188156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188156));
	wire w192156;
	repeater #(2, 1'b0, 0, 0) c192156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192156));
	wire w196156;
	repeater #(2, 1'b0, 0, 0) c196156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196156));
	wire w37158;
	repeater #(1, 1'b0, 0, 0) c37158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37158));
	wire w39158;
	torch #(1'b0) c39158 (.i_clk(tick), .i_in(), .o_out(w39158));
	wire w45158;
	torch #(1'b1) c45158 (.i_clk(tick), .i_in(), .o_out(w45158));
	wire w53158;
	repeater #(1, 1'b0, 0, 0) c53158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53158));
	wire w55158;
	torch #(1'b0) c55158 (.i_clk(tick), .i_in(), .o_out(w55158));
	wire w71158;
	repeater #(1, 1'b0, 0, 0) c71158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71158));
	wire w73158;
	torch #(1'b0) c73158 (.i_clk(tick), .i_in(), .o_out(w73158));
	wire w79158;
	torch #(1'b1) c79158 (.i_clk(tick), .i_in(), .o_out(w79158));
	wire w87158;
	repeater #(1, 1'b0, 0, 0) c87158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87158));
	wire w89158;
	torch #(1'b0) c89158 (.i_clk(tick), .i_in(), .o_out(w89158));
	wire w41160;
	repeater #(1, 1'b0, 0, 0) c41160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41160));
	wire w57160;
	repeater #(1, 1'b0, 0, 0) c57160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57160));
	wire w75160;
	repeater #(1, 1'b0, 0, 0) c75160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75160));
	wire w91160;
	repeater #(1, 1'b0, 0, 0) c91160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91160));
	wire w38162;
	torch #(1'b1) c38162 (.i_clk(tick), .i_in(), .o_out(w38162));
	wire w54162;
	torch #(1'b1) c54162 (.i_clk(tick), .i_in(), .o_out(w54162));
	wire w72162;
	torch #(1'b1) c72162 (.i_clk(tick), .i_in(), .o_out(w72162));
	wire w88162;
	torch #(1'b1) c88162 (.i_clk(tick), .i_in(), .o_out(w88162));
	wire w46164;
	torch #(1'b1) c46164 (.i_clk(tick), .i_in(), .o_out(w46164));
	wire w80164;
	torch #(1'b1) c80164 (.i_clk(tick), .i_in(), .o_out(w80164));
	wire w37165;
	repeater #(1, 1'b0, 0, 0) c37165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37165));
	wire w49165;
	repeater #(1, 1'b0, 0, 0) c49165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49165));
	wire w71165;
	repeater #(1, 1'b0, 0, 0) c71165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71165));
	wire w83165;
	repeater #(1, 1'b0, 0, 0) c83165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83165));
	wire w43166;
	repeater #(1, 1'b0, 0, 0) c43166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43166));
	wire w77166;
	repeater #(1, 1'b0, 0, 0) c77166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77166));
	wire w43168;
	repeater #(1, 1'b0, 0, 0) c43168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43168));
	wire w77168;
	repeater #(1, 1'b0, 0, 0) c77168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77168));
	wire w131106;
	repeater #(1, 1'b0, 0, 0) c131106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131106));
	wire w131122;
	repeater #(1, 1'b0, 0, 0) c131122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131122));
	wire w11126;
	repeater #(1, 1'b0, 0, 0) c11126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11126));
	wire w1681135;
	repeater #(1, 1'b0, 0, 0) c1681135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1681135));
	wire w1721135;
	repeater #(1, 1'b0, 0, 0) c1721135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1721135));
	wire w1761135;
	repeater #(1, 1'b0, 0, 0) c1761135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1761135));
	wire w1801135;
	repeater #(1, 1'b0, 0, 0) c1801135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1801135));
	wire w1841135;
	repeater #(1, 1'b0, 0, 0) c1841135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1841135));
	wire w1881135;
	repeater #(1, 1'b0, 0, 0) c1881135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1881135));
	wire w1921135;
	repeater #(1, 1'b0, 0, 0) c1921135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1921135));
	wire w178047;

	wire w176049;

	wire w174051;

	wire w172053;

	wire w170055;

	wire w28060;
	repeater #(2, 1'b0, 0, 0) c28060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28060));
	wire w62060;
	repeater #(2, 1'b0, 0, 0) c62060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62060));
	wire w20062;
	torch #(1'b1) c20062 (.i_clk(tick), .i_in(), .o_out(w20062));
	wire w30062;
	repeater #(1, 1'b0, 0, 0) c30062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30062));
	wire w36062;
	torch #(1'b1) c36062 (.i_clk(tick), .i_in(), .o_out(w36062));
	wire w54062;
	torch #(1'b1) c54062 (.i_clk(tick), .i_in(), .o_out(w54062));
	wire w64062;
	repeater #(1, 1'b1, 0, 0) c64062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64062));
	wire w70062;
	torch #(1'b1) c70062 (.i_clk(tick), .i_in(), .o_out(w70062));
	wire w30066;
	repeater #(1, 1'b0, 0, 0) c30066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30066));
	wire w64066;
	repeater #(1, 1'b1, 0, 0) c64066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64066));
	wire w19067;

	wire w35067;

	wire w53067;

	wire w69067;

	wire w27068;

	wire w61068;

	wire w24069;

	wire w29069;

	wire w30069;

	wire w58069;

	wire w63069;

	wire w64069;

	wire w19070;

	wire w53070;

	wire w156070;
	repeater #(1, 1'b0, 0, 0) c156070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156070));
	wire w176070;
	repeater #(1, 1'b0, 0, 0) c176070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176070));
	wire w22071;

	wire w38071;

	wire w56071;

	wire w72071;

	wire w28072;

	wire w29072;

	wire w62072;

	wire w63072;

	wire w14073;

	wire w48073;

	wire w15075;
	repeater #(1, 1'b1, 0, 0) c15075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15075));
	wire w19075;
	repeater #(1, 1'b1, 0, 0) c19075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19075));
	wire w23075;
	repeater #(1, 1'b1, 0, 0) c23075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23075));
	wire w27075;
	repeater #(1, 1'b0, 0, 0) c27075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27075));
	wire w31075;
	repeater #(1, 1'b1, 0, 0) c31075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31075));
	wire w35075;
	repeater #(1, 1'b1, 0, 0) c35075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35075));
	wire w39075;
	repeater #(1, 1'b1, 0, 0) c39075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39075));
	wire w49075;
	repeater #(1, 1'b1, 0, 0) c49075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49075));
	wire w53075;
	repeater #(1, 1'b1, 0, 0) c53075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53075));
	wire w57075;
	repeater #(1, 1'b0, 0, 0) c57075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57075));
	wire w61075;
	repeater #(1, 1'b1, 0, 0) c61075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61075));
	wire w65075;
	repeater #(1, 1'b0, 0, 0) c65075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65075));
	wire w69075;
	repeater #(1, 1'b1, 0, 0) c69075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69075));
	wire w73075;
	repeater #(1, 1'b1, 0, 0) c73075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73075));
	wire w22084;

	wire w56084;

	wire w20085;
	repeater #(1, 1'b1, 0, 0) c20085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20085));
	wire w36085;
	repeater #(1, 1'b1, 0, 0) c36085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36085));
	wire w54085;
	repeater #(1, 1'b1, 0, 0) c54085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54085));
	wire w70085;
	repeater #(1, 1'b1, 0, 0) c70085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70085));
	wire w11086;
	repeater #(1, 1'b1, 0, 0) c11086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11086));
	wire w27086;
	repeater #(1, 1'b1, 0, 0) c27086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27086));
	wire w45086;
	repeater #(1, 1'b1, 0, 0) c45086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45086));
	wire w61086;
	repeater #(1, 1'b0, 0, 0) c61086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61086));
	wire w156086;
	repeater #(1, 1'b0, 0, 0) c156086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156086));
	wire w176086;
	repeater #(1, 1'b0, 0, 0) c176086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176086));
	wire w22087;

	wire w38087;

	wire w56087;

	wire w72087;

	wire w30088;

	wire w64088;

	wire w11089;

	wire w25089;

	wire w27089;

	wire w28089;

	wire w33089;

	wire w41089;

	wire w45089;

	wire w59089;

	wire w61089;

	wire w62089;

	wire w67089;

	wire w75089;

	wire w38090;

	wire w72090;

	wire w19091;

	wire w35091;

	wire w36091;

	wire w53091;

	wire w69091;

	wire w70091;

	wire w11093;

	wire w12093;

	wire w25093;

	wire w27093;

	wire w28093;

	wire w41093;

	wire w45093;

	wire w46093;

	wire w59093;

	wire w61093;

	wire w62093;

	wire w75093;

	wire w22095;
	torch #(1'b1) c22095 (.i_clk(tick), .i_in(), .o_out(w22095));
	wire w23095;

	wire w28095;

	wire w56095;
	torch #(1'b1) c56095 (.i_clk(tick), .i_in(), .o_out(w56095));
	wire w57095;

	wire w62095;

	wire w23096;

	wire w25096;

	wire w39096;

	wire w41096;

	wire w57096;

	wire w59096;

	wire w73096;

	wire w75096;

	wire w25098;

	wire w26098;

	wire w27098;

	wire w41098;

	wire w42098;

	wire w43098;

	wire w59098;

	wire w60098;

	wire w61098;

	wire w75098;

	wire w76098;

	wire w77098;

	wire w20099;

	wire w21099;

	wire w27099;

	wire w36099;

	wire w37099;

	wire w43099;

	wire w54099;

	wire w55099;

	wire w61099;

	wire w70099;

	wire w71099;

	wire w77099;

	wire w170101;
	torch #(1'b0) c170101 (.i_clk(tick), .i_in(), .o_out(w170101));
	wire w250101;
	repeater #(1, 1'b0, 0, 0) c250101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250101));
	wire w270101;
	torch #(1'b0) c270101 (.i_clk(tick), .i_in(), .o_out(w270101));
	wire w330101;
	torch #(1'b1) c330101 (.i_clk(tick), .i_in(), .o_out(w330101));
	wire w410101;
	repeater #(1, 1'b0, 0, 0) c410101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w410101));
	wire w430101;
	torch #(1'b0) c430101 (.i_clk(tick), .i_in(), .o_out(w430101));
	wire w510101;
	torch #(1'b0) c510101 (.i_clk(tick), .i_in(), .o_out(w510101));
	wire w590101;
	repeater #(1, 1'b0, 0, 0) c590101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590101));
	wire w610101;
	torch #(1'b0) c610101 (.i_clk(tick), .i_in(), .o_out(w610101));
	wire w670101;
	torch #(1'b1) c670101 (.i_clk(tick), .i_in(), .o_out(w670101));
	wire w750101;
	repeater #(1, 1'b0, 0, 0) c750101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w750101));
	wire w770101;
	torch #(1'b0) c770101 (.i_clk(tick), .i_in(), .o_out(w770101));
	wire w1560102;
	repeater #(1, 1'b0, 0, 0) c1560102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560102));
	wire w1760102;
	repeater #(1, 1'b0, 0, 0) c1760102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1760102));
	wire w290103;
	repeater #(1, 1'b1, 0, 0) c290103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290103));
	wire w630103;
	repeater #(1, 1'b1, 0, 0) c630103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630103));
	wire w260105;
	torch #(1'b1) c260105 (.i_clk(tick), .i_in(), .o_out(w260105));
	wire w420105;
	torch #(1'b1) c420105 (.i_clk(tick), .i_in(), .o_out(w420105));
	wire w600105;
	torch #(1'b1) c600105 (.i_clk(tick), .i_in(), .o_out(w600105));
	wire w760105;
	torch #(1'b1) c760105 (.i_clk(tick), .i_in(), .o_out(w760105));
	wire w180107;
	torch #(1'b1) c180107 (.i_clk(tick), .i_in(), .o_out(w180107));
	wire w340107;
	torch #(1'b1) c340107 (.i_clk(tick), .i_in(), .o_out(w340107));
	wire w520107;
	torch #(1'b1) c520107 (.i_clk(tick), .i_in(), .o_out(w520107));
	wire w680107;
	torch #(1'b1) c680107 (.i_clk(tick), .i_in(), .o_out(w680107));
	wire w250108;
	repeater #(1, 1'b0, 0, 0) c250108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250108));
	wire w370108;
	repeater #(1, 1'b0, 0, 0) c370108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370108));
	wire w590108;
	repeater #(1, 1'b0, 0, 0) c590108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590108));
	wire w710108;
	repeater #(1, 1'b0, 0, 0) c710108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710108));
	wire w190109;
	repeater #(1, 1'b0, 0, 0) c190109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190109));
	wire w310109;
	repeater #(1, 1'b0, 0, 0) c310109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310109));
	wire w530109;
	repeater #(1, 1'b0, 0, 0) c530109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530109));
	wire w650109;
	repeater #(1, 1'b0, 0, 0) c650109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650109));
	wire w310111;
	repeater #(1, 1'b0, 0, 0) c310111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310111));
	wire w650111;
	repeater #(1, 1'b0, 0, 0) c650111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650111));
	wire w1560118;
	repeater #(1, 1'b0, 0, 0) c1560118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560118));
	wire w1760118;
	repeater #(1, 1'b0, 0, 0) c1760118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1760118));
	wire w1560134;
	repeater #(1, 1'b0, 0, 0) c1560134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560134));
	wire w1760134;
	repeater #(1, 1'b0, 0, 0) c1760134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1760134));
	wire w1880159;
	torch #(1'b1) c1880159 (.i_clk(tick), .i_in(), .o_out(w1880159));
	wire w1820163;
	torch #(1'b1) c1820163 (.i_clk(tick), .i_in(), .o_out(w1820163));
	wire w156111;
	repeater #(1, 1'b0, 0, 0) c156111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156111));
	wire w160111;
	repeater #(1, 1'b0, 0, 0) c160111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160111));
	wire w164111;
	repeater #(1, 1'b0, 0, 0) c164111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164111));
	wire w168111;
	repeater #(1, 1'b0, 0, 0) c168111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168111));
	wire w172111;
	repeater #(1, 1'b0, 0, 0) c172111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172111));
	wire w176111;
	repeater #(1, 1'b0, 0, 0) c176111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176111));
	wire w180111;
	repeater #(1, 1'b0, 0, 0) c180111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180111));
	wire w153121;
	repeater #(1, 1'b0, 0, 0) c153121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153121));
	wire w157121;
	repeater #(1, 1'b0, 0, 0) c157121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157121));
	wire w161121;
	repeater #(1, 1'b1, 0, 0) c161121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161121));
	wire w165121;
	repeater #(1, 1'b0, 0, 0) c165121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165121));
	wire w169121;
	repeater #(1, 1'b1, 0, 0) c169121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169121));
	wire w173121;
	repeater #(1, 1'b0, 0, 0) c173121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173121));
	wire w177121;
	repeater #(1, 1'b0, 0, 0) c177121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177121));
	wire w153124;
	torch #(1'b1) c153124 (.i_clk(tick), .i_in(), .o_out(w153124));
	wire w157124;
	torch #(1'b1) c157124 (.i_clk(tick), .i_in(), .o_out(w157124));
	wire w161124;
	torch #(1'b0) c161124 (.i_clk(tick), .i_in(), .o_out(w161124));
	wire w165124;
	torch #(1'b1) c165124 (.i_clk(tick), .i_in(), .o_out(w165124));
	wire w169124;
	torch #(1'b0) c169124 (.i_clk(tick), .i_in(), .o_out(w169124));
	wire w173124;
	torch #(1'b1) c173124 (.i_clk(tick), .i_in(), .o_out(w173124));
	wire w177124;
	torch #(1'b1) c177124 (.i_clk(tick), .i_in(), .o_out(w177124));
	wire w164127;
	repeater #(1, 1'b0, 0, 0) c164127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164127));
	wire w166127;
	repeater #(1, 1'b1, 0, 0) c166127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166127));
	wire w168127;
	repeater #(1, 1'b0, 0, 0) c168127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168127));
	wire w170127;
	repeater #(1, 1'b0, 0, 0) c170127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170127));
	wire w172127;
	repeater #(1, 1'b1, 0, 0) c172127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172127));
	wire w174127;
	repeater #(1, 1'b1, 0, 0) c174127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174127));
	wire w176127;
	repeater #(1, 1'b1, 0, 0) c176127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176127));
	wire w178127;
	repeater #(1, 1'b1, 0, 0) c178127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178127));
	wire w162129;
	repeater #(1, 1'b0, 0, 0) c162129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162129));
	wire w160131;
	repeater #(1, 1'b0, 0, 0) c160131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160131));
	wire w158133;
	repeater #(1, 1'b1, 0, 0) c158133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158133));
	wire w156135;
	repeater #(1, 1'b1, 0, 0) c156135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156135));
	wire w154137;
	repeater #(1, 1'b1, 0, 0) c154137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154137));
	wire w152139;
	repeater #(1, 1'b1, 0, 0) c152139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152139));
	wire w42145;
	torch #(1'b1) c42145 (.i_clk(tick), .i_in(), .o_out(w42145));
	wire w76145;
	repeater #(1, 1'b1, 0, 0) c76145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76145));
	wire w110145;
	torch #(1'b1) c110145 (.i_clk(tick), .i_in(), .o_out(w110145));
	wire w144145;
	repeater #(1, 1'b1, 0, 0) c144145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144145));
	wire w40147;
	repeater #(1, 1'b1, 0, 0) c40147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40147));
	wire w74147;
	repeater #(1, 1'b1, 0, 0) c74147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74147));
	wire w108147;
	repeater #(1, 1'b1, 0, 0) c108147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108147));
	wire w142147;
	repeater #(1, 1'b1, 0, 0) c142147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142147));
	wire w178148;
	repeater #(1, 1'b1, 0, 0) c178148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178148));
	wire w38149;
	torch #(1'b1) c38149 (.i_clk(tick), .i_in(), .o_out(w38149));
	wire w72149;
	repeater #(1, 1'b1, 0, 0) c72149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72149));
	wire w106149;
	torch #(1'b1) c106149 (.i_clk(tick), .i_in(), .o_out(w106149));
	wire w140149;
	repeater #(1, 1'b1, 0, 0) c140149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140149));
	wire w176150;
	repeater #(1, 1'b1, 0, 0) c176150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176150));
	wire w36151;
	repeater #(1, 1'b1, 0, 0) c36151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36151));
	wire w70151;
	repeater #(1, 1'b1, 0, 0) c70151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70151));
	wire w104151;
	repeater #(1, 1'b1, 0, 0) c104151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104151));
	wire w138151;
	repeater #(1, 1'b1, 0, 0) c138151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138151));
	wire w184151;
	repeater #(1, 1'b1, 0, 0) c184151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184151));
	wire w174152;
	repeater #(1, 1'b1, 0, 0) c174152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174152));
	wire w34153;
	torch #(1'b0) c34153 (.i_clk(tick), .i_in(), .o_out(w34153));
	wire w68153;
	repeater #(1, 1'b0, 0, 0) c68153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68153));
	wire w102153;
	torch #(1'b0) c102153 (.i_clk(tick), .i_in(), .o_out(w102153));
	wire w136153;
	repeater #(1, 1'b0, 0, 0) c136153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136153));
	wire w172154;
	repeater #(1, 1'b1, 0, 0) c172154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172154));
	wire w32155;
	repeater #(1, 1'b0, 0, 0) c32155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32155));
	wire w66155;
	repeater #(1, 1'b0, 0, 0) c66155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66155));
	wire w100155;
	repeater #(1, 1'b0, 0, 0) c100155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100155));
	wire w134155;
	repeater #(1, 1'b0, 0, 0) c134155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134155));
	wire w16156;
	repeater #(1, 1'b1, 0, 0) c16156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16156));
	wire w18156;
	torch #(1'b1) c18156 (.i_clk(tick), .i_in(), .o_out(w18156));
	wire w20156;
	repeater #(1, 1'b1, 0, 0) c20156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20156));
	wire w22156;
	torch #(1'b1) c22156 (.i_clk(tick), .i_in(), .o_out(w22156));
	wire w24156;
	repeater #(1, 1'b0, 0, 0) c24156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24156));
	wire w26156;
	torch #(1'b0) c26156 (.i_clk(tick), .i_in(), .o_out(w26156));
	wire w28156;
	repeater #(1, 1'b0, 0, 0) c28156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28156));
	wire w30156;
	torch #(1'b1) c30156 (.i_clk(tick), .i_in(), .o_out(w30156));
	wire w50156;
	repeater #(1, 1'b1, 0, 0) c50156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50156));
	wire w52156;
	repeater #(1, 1'b1, 0, 0) c52156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52156));
	wire w54156;
	repeater #(1, 1'b1, 0, 0) c54156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54156));
	wire w56156;
	repeater #(1, 1'b1, 0, 0) c56156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56156));
	wire w58156;
	repeater #(1, 1'b0, 0, 0) c58156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58156));
	wire w60156;
	repeater #(1, 1'b0, 0, 0) c60156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60156));
	wire w62156;
	repeater #(1, 1'b0, 0, 0) c62156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62156));
	wire w64156;
	repeater #(1, 1'b1, 0, 0) c64156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64156));
	wire w86156;
	torch #(1'b1) c86156 (.i_clk(tick), .i_in(), .o_out(w86156));
	wire w90156;
	torch #(1'b1) c90156 (.i_clk(tick), .i_in(), .o_out(w90156));
	wire w94156;
	torch #(1'b0) c94156 (.i_clk(tick), .i_in(), .o_out(w94156));
	wire w98156;
	torch #(1'b1) c98156 (.i_clk(tick), .i_in(), .o_out(w98156));
	wire w118156;
	repeater #(1, 1'b1, 0, 0) c118156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118156));
	wire w120156;
	repeater #(1, 1'b1, 0, 0) c120156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120156));
	wire w122156;
	repeater #(1, 1'b1, 0, 0) c122156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122156));
	wire w124156;
	repeater #(1, 1'b1, 0, 0) c124156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124156));
	wire w126156;
	repeater #(1, 1'b0, 0, 0) c126156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126156));
	wire w128156;
	repeater #(1, 1'b0, 0, 0) c128156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128156));
	wire w130156;
	repeater #(1, 1'b0, 0, 0) c130156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130156));
	wire w132156;
	repeater #(1, 1'b1, 0, 0) c132156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132156));
	wire w170156;
	repeater #(1, 1'b0, 0, 0) c170156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170156));
	wire w85157;
	repeater #(1, 1'b1, 0, 0) c85157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85157));
	wire w89157;
	repeater #(1, 1'b1, 0, 0) c89157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89157));
	wire w93157;
	repeater #(1, 1'b0, 0, 0) c93157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93157));
	wire w97157;
	repeater #(1, 1'b0, 0, 0) c97157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97157));
	wire w156157;
	repeater #(1, 1'b1, 0, 0) c156157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156157));
	wire w158157;
	repeater #(1, 1'b1, 0, 0) c158157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158157));
	wire w160157;
	repeater #(1, 1'b0, 0, 0) c160157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160157));
	wire w162157;
	repeater #(1, 1'b0, 0, 0) c162157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162157));
	wire w164157;
	repeater #(1, 1'b0, 0, 0) c164157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164157));
	wire w166157;
	repeater #(1, 1'b1, 0, 0) c166157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166157));
	wire w168157;
	repeater #(1, 1'b0, 0, 0) c168157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168157));
	wire w86159;
	torch #(1'b1) c86159 (.i_clk(tick), .i_in(), .o_out(w86159));
	wire w90159;
	torch #(1'b1) c90159 (.i_clk(tick), .i_in(), .o_out(w90159));
	wire w94159;
	torch #(1'b1) c94159 (.i_clk(tick), .i_in(), .o_out(w94159));
	wire w98159;
	torch #(1'b0) c98159 (.i_clk(tick), .i_in(), .o_out(w98159));
	wire w102159;
	torch #(1'b1) c102159 (.i_clk(tick), .i_in(), .o_out(w102159));
	wire w106159;
	torch #(1'b1) c106159 (.i_clk(tick), .i_in(), .o_out(w106159));
	wire w110159;
	torch #(1'b1) c110159 (.i_clk(tick), .i_in(), .o_out(w110159));
	wire w120159;
	torch #(1'b1) c120159 (.i_clk(tick), .i_in(), .o_out(w120159));
	wire w124159;
	torch #(1'b1) c124159 (.i_clk(tick), .i_in(), .o_out(w124159));
	wire w128159;
	torch #(1'b0) c128159 (.i_clk(tick), .i_in(), .o_out(w128159));
	wire w132159;
	torch #(1'b1) c132159 (.i_clk(tick), .i_in(), .o_out(w132159));
	wire w136159;
	torch #(1'b0) c136159 (.i_clk(tick), .i_in(), .o_out(w136159));
	wire w140159;
	torch #(1'b1) c140159 (.i_clk(tick), .i_in(), .o_out(w140159));
	wire w144159;
	torch #(1'b1) c144159 (.i_clk(tick), .i_in(), .o_out(w144159));
	wire w16160;
	repeater #(2, 1'b1, 0, 0) c16160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16160));
	wire w20160;
	repeater #(2, 1'b1, 0, 0) c20160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20160));
	wire w24160;
	repeater #(2, 1'b0, 0, 0) c24160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24160));
	wire w40160;
	repeater #(2, 1'b1, 0, 0) c40160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40160));
	wire w50160;
	repeater #(2, 1'b1, 0, 0) c50160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50160));
	wire w54160;
	repeater #(2, 1'b1, 0, 0) c54160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54160));
	wire w58160;
	repeater #(2, 1'b0, 0, 0) c58160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58160));
	wire w74160;
	repeater #(2, 1'b1, 0, 0) c74160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74160));
	wire w16162;
	torch #(1'b1) c16162 (.i_clk(tick), .i_in(), .o_out(w16162));
	wire w26162;
	repeater #(1, 1'b1, 0, 0) c26162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26162));
	wire w32162;
	torch #(1'b1) c32162 (.i_clk(tick), .i_in(), .o_out(w32162));
	wire w42162;
	repeater #(1, 1'b1, 0, 0) c42162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42162));
	wire w50162;
	torch #(1'b1) c50162 (.i_clk(tick), .i_in(), .o_out(w50162));
	wire w60162;
	repeater #(1, 1'b0, 0, 0) c60162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60162));
	wire w66162;
	torch #(1'b1) c66162 (.i_clk(tick), .i_in(), .o_out(w66162));
	wire w76162;
	repeater #(1, 1'b1, 0, 0) c76162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76162));
	wire w91163;
	torch #(1'b1) c91163 (.i_clk(tick), .i_in(), .o_out(w91163));
	wire w95163;
	torch #(1'b1) c95163 (.i_clk(tick), .i_in(), .o_out(w95163));
	wire w99163;
	torch #(1'b1) c99163 (.i_clk(tick), .i_in(), .o_out(w99163));
	wire w103163;
	torch #(1'b1) c103163 (.i_clk(tick), .i_in(), .o_out(w103163));
	wire w127163;
	torch #(1'b1) c127163 (.i_clk(tick), .i_in(), .o_out(w127163));
	wire w131163;
	torch #(1'b1) c131163 (.i_clk(tick), .i_in(), .o_out(w131163));
	wire w135163;
	torch #(1'b1) c135163 (.i_clk(tick), .i_in(), .o_out(w135163));
	wire w139163;
	torch #(1'b1) c139163 (.i_clk(tick), .i_in(), .o_out(w139163));
	wire w17165;
	repeater #(1, 1'b1, 0, 0) c17165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17165));
	wire w33165;
	repeater #(1, 1'b1, 0, 0) c33165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33165));
	wire w51165;
	repeater #(1, 1'b1, 0, 0) c51165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51165));
	wire w67165;
	repeater #(1, 1'b1, 0, 0) c67165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67165));
	wire w26166;
	repeater #(1, 1'b1, 0, 0) c26166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26166));
	wire w42166;
	repeater #(1, 1'b1, 0, 0) c42166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42166));
	wire w60166;
	repeater #(1, 1'b0, 0, 0) c60166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60166));
	wire w76166;
	repeater #(1, 1'b1, 0, 0) c76166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76166));
	wire w15167;

	wire w31167;

	wire w49167;

	wire w65167;

	wire w154167;
	repeater #(1, 1'b1, 0, 0) c154167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154167));
	wire w158167;
	repeater #(1, 1'b1, 0, 0) c158167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158167));
	wire w162167;
	repeater #(1, 1'b1, 0, 0) c162167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162167));
	wire w166167;
	repeater #(1, 1'b0, 0, 0) c166167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166167));
	wire w170167;
	repeater #(1, 1'b1, 0, 0) c170167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170167));
	wire w174167;
	repeater #(1, 1'b1, 0, 0) c174167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174167));
	wire w178167;
	repeater #(1, 1'b1, 0, 0) c178167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178167));
	wire w23168;

	wire w57168;

	wire w20169;

	wire w25169;

	wire w26169;

	wire w42169;

	wire w54169;

	wire w59169;

	wire w60169;

	wire w76169;

	wire w184169;
	repeater #(1, 1'b1, 0, 0) c184169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184169));
	wire w15170;

	wire w49170;

	wire w18171;

	wire w34171;

	wire w52171;

	wire w68171;

	wire w181171;
	repeater #(1, 1'b0, 0, 0) c181171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181171));
	wire w24172;

	wire w25172;

	wire w40172;

	wire w41172;

	wire w58172;

	wire w59172;

	wire w74172;

	wire w75172;

	wire w34173;

	wire w38173;

	wire w68173;

	wire w72173;

	wire w151173;
	repeater #(1, 1'b0, 0, 0) c151173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151173));
	wire w160176;
	torch #(1'b1) c160176 (.i_clk(tick), .i_in(), .o_out(w160176));
	wire w164176;
	torch #(1'b1) c164176 (.i_clk(tick), .i_in(), .o_out(w164176));
	wire w168176;
	torch #(1'b1) c168176 (.i_clk(tick), .i_in(), .o_out(w168176));
	wire w172176;
	torch #(1'b1) c172176 (.i_clk(tick), .i_in(), .o_out(w172176));
	wire w15177;

	wire w16177;

	wire w19177;

	wire w20177;

	wire w23177;

	wire w24177;

	wire w27177;

	wire w28177;

	wire w31177;

	wire w32177;

	wire w35177;

	wire w36177;

	wire w39177;

	wire w40177;

	wire w49177;

	wire w50177;

	wire w53177;

	wire w54177;

	wire w57177;

	wire w58177;

	wire w61177;

	wire w62177;

	wire w65177;

	wire w66177;

	wire w69177;

	wire w70177;

	wire w73177;

	wire w74177;

	wire w16179;

	wire w20179;

	wire w24179;

	wire w28179;

	wire w32179;

	wire w36179;

	wire w40179;

	wire w50179;

	wire w54179;

	wire w58179;

	wire w62179;

	wire w66179;

	wire w70179;

	wire w74179;

	wire w153180;
	torch #(1'b0) c153180 (.i_clk(tick), .i_in(), .o_out(w153180));
	wire w157180;
	torch #(1'b0) c157180 (.i_clk(tick), .i_in(), .o_out(w157180));
	wire w161180;
	torch #(1'b0) c161180 (.i_clk(tick), .i_in(), .o_out(w161180));
	wire w165180;
	torch #(1'b1) c165180 (.i_clk(tick), .i_in(), .o_out(w165180));
	wire w169180;
	torch #(1'b0) c169180 (.i_clk(tick), .i_in(), .o_out(w169180));
	wire w173180;
	torch #(1'b0) c173180 (.i_clk(tick), .i_in(), .o_out(w173180));
	wire w177180;
	torch #(1'b0) c177180 (.i_clk(tick), .i_in(), .o_out(w177180));
	wire w14182;

	wire w18182;

	wire w22182;

	wire w26182;

	wire w48182;

	wire w52182;

	wire w56182;

	wire w60182;

	wire w154182;
	torch #(1'b1) c154182 (.i_clk(tick), .i_in(), .o_out(w154182));
	wire w158182;
	torch #(1'b1) c158182 (.i_clk(tick), .i_in(), .o_out(w158182));
	wire w162182;
	torch #(1'b1) c162182 (.i_clk(tick), .i_in(), .o_out(w162182));
	wire w166182;
	torch #(1'b1) c166182 (.i_clk(tick), .i_in(), .o_out(w166182));
	wire w170182;
	torch #(1'b1) c170182 (.i_clk(tick), .i_in(), .o_out(w170182));
	wire w174182;
	torch #(1'b1) c174182 (.i_clk(tick), .i_in(), .o_out(w174182));
	wire w178182;
	torch #(1'b1) c178182 (.i_clk(tick), .i_in(), .o_out(w178182));
	wire w26184;

	wire w60184;

	wire w155184;
	torch #(1'b0) c155184 (.i_clk(tick), .i_in(), .o_out(w155184));
	wire w159184;
	torch #(1'b0) c159184 (.i_clk(tick), .i_in(), .o_out(w159184));
	wire w163184;
	torch #(1'b0) c163184 (.i_clk(tick), .i_in(), .o_out(w163184));
	wire w167184;
	torch #(1'b0) c167184 (.i_clk(tick), .i_in(), .o_out(w167184));
	wire w171184;
	torch #(1'b0) c171184 (.i_clk(tick), .i_in(), .o_out(w171184));
	wire w175184;
	torch #(1'b0) c175184 (.i_clk(tick), .i_in(), .o_out(w175184));
	wire w179184;
	torch #(1'b0) c179184 (.i_clk(tick), .i_in(), .o_out(w179184));
	wire w24185;
	repeater #(1, 1'b1, 0, 0) c24185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24185));
	wire w58185;
	repeater #(1, 1'b0, 0, 0) c58185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58185));
	wire w15186;
	repeater #(1, 1'b1, 0, 0) c15186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15186));
	wire w31186;
	repeater #(1, 1'b1, 0, 0) c31186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31186));
	wire w49186;
	repeater #(1, 1'b1, 0, 0) c49186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49186));
	wire w65186;
	repeater #(1, 1'b1, 0, 0) c65186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65186));
	wire w186186;
	repeater #(1, 1'b1, 0, 0) c186186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186186));
	wire w188186;
	repeater #(1, 1'b1, 0, 0) c188186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188186));
	wire w190186;
	repeater #(1, 1'b1, 0, 0) c190186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190186));
	wire w26187;

	wire w60187;

	wire w181187;
	repeater #(1, 1'b0, 0, 0) c181187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181187));
	wire w184187;
	repeater #(1, 1'b1, 0, 0) c184187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184187));
	wire w18188;

	wire w34188;

	wire w52188;

	wire w68188;

	wire w15189;

	wire w21189;

	wire w29189;

	wire w31189;

	wire w32189;

	wire w37189;

	wire w49189;

	wire w55189;

	wire w63189;

	wire w65189;

	wire w66189;

	wire w71189;

	wire w151189;
	repeater #(1, 1'b0, 0, 0) c151189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151189));
	wire w23191;

	wire w24191;

	wire w39191;

	wire w40191;

	wire w57191;

	wire w58191;

	wire w73191;

	wire w74191;

	wire w160192;
	torch #(1'b1) c160192 (.i_clk(tick), .i_in(), .o_out(w160192));
	wire w164192;
	torch #(1'b1) c164192 (.i_clk(tick), .i_in(), .o_out(w164192));
	wire w168192;
	torch #(1'b1) c168192 (.i_clk(tick), .i_in(), .o_out(w168192));
	wire w172192;
	torch #(1'b1) c172192 (.i_clk(tick), .i_in(), .o_out(w172192));
	wire w15193;

	wire w16193;

	wire w29193;

	wire w31193;

	wire w32193;

	wire w49193;

	wire w50193;

	wire w63193;

	wire w65193;

	wire w66193;

	wire w26195;
	torch #(1'b1) c26195 (.i_clk(tick), .i_in(), .o_out(w26195));
	wire w27195;

	wire w32195;

	wire w60195;
	torch #(1'b1) c60195 (.i_clk(tick), .i_in(), .o_out(w60195));
	wire w61195;

	wire w66195;

	wire w27196;

	wire w29196;

	wire w61196;

	wire w63196;

	wire w153196;
	torch #(1'b0) c153196 (.i_clk(tick), .i_in(), .o_out(w153196));
	wire w157196;
	torch #(1'b0) c157196 (.i_clk(tick), .i_in(), .o_out(w157196));
	wire w161196;
	torch #(1'b1) c161196 (.i_clk(tick), .i_in(), .o_out(w161196));
	wire w165196;
	torch #(1'b0) c165196 (.i_clk(tick), .i_in(), .o_out(w165196));
	wire w169196;
	torch #(1'b1) c169196 (.i_clk(tick), .i_in(), .o_out(w169196));
	wire w173196;
	torch #(1'b0) c173196 (.i_clk(tick), .i_in(), .o_out(w173196));
	wire w177196;
	torch #(1'b0) c177196 (.i_clk(tick), .i_in(), .o_out(w177196));
	wire w29198;

	wire w30198;

	wire w31198;

	wire w63198;

	wire w64198;

	wire w65198;

	wire w99198;
	repeater #(1, 1'b0, 0, 0) c99198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99198));
	wire w131198;
	repeater #(1, 1'b0, 0, 0) c131198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131198));
	wire w154198;
	torch #(1'b1) c154198 (.i_clk(tick), .i_in(), .o_out(w154198));
	wire w158198;
	torch #(1'b1) c158198 (.i_clk(tick), .i_in(), .o_out(w158198));
	wire w162198;
	torch #(1'b1) c162198 (.i_clk(tick), .i_in(), .o_out(w162198));
	wire w166198;
	torch #(1'b1) c166198 (.i_clk(tick), .i_in(), .o_out(w166198));
	wire w170198;
	torch #(1'b1) c170198 (.i_clk(tick), .i_in(), .o_out(w170198));
	wire w174198;
	torch #(1'b1) c174198 (.i_clk(tick), .i_in(), .o_out(w174198));
	wire w178198;
	torch #(1'b1) c178198 (.i_clk(tick), .i_in(), .o_out(w178198));
	wire w24199;

	wire w25199;

	wire w31199;

	wire w40199;

	wire w41199;

	wire w58199;

	wire w59199;

	wire w65199;

	wire w74199;

	wire w75199;

	wire w96199;

	wire w134199;

	wire w951100;
	repeater #(2, 1'b0, 0, 0) c951100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951100));
	wire w1351100;
	repeater #(2, 1'b0, 0, 0) c1351100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1351100));
	wire w1551100;
	torch #(1'b0) c1551100 (.i_clk(tick), .i_in(), .o_out(w1551100));
	wire w1591100;
	torch #(1'b0) c1591100 (.i_clk(tick), .i_in(), .o_out(w1591100));
	wire w1631100;
	torch #(1'b0) c1631100 (.i_clk(tick), .i_in(), .o_out(w1631100));
	wire w1671100;
	torch #(1'b0) c1671100 (.i_clk(tick), .i_in(), .o_out(w1671100));
	wire w1711100;
	torch #(1'b0) c1711100 (.i_clk(tick), .i_in(), .o_out(w1711100));
	wire w1751100;
	torch #(1'b0) c1751100 (.i_clk(tick), .i_in(), .o_out(w1751100));
	wire w1791100;
	torch #(1'b0) c1791100 (.i_clk(tick), .i_in(), .o_out(w1791100));
	wire w211101;
	torch #(1'b0) c211101 (.i_clk(tick), .i_in(), .o_out(w211101));
	wire w291101;
	repeater #(1, 1'b1, 0, 0) c291101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w291101));
	wire w311101;
	torch #(1'b0) c311101 (.i_clk(tick), .i_in(), .o_out(w311101));
	wire w371101;
	torch #(1'b0) c371101 (.i_clk(tick), .i_in(), .o_out(w371101));
	wire w551101;
	torch #(1'b0) c551101 (.i_clk(tick), .i_in(), .o_out(w551101));
	wire w631101;
	repeater #(1, 1'b1, 0, 0) c631101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w631101));
	wire w651101;
	torch #(1'b0) c651101 (.i_clk(tick), .i_in(), .o_out(w651101));
	wire w711101;
	torch #(1'b0) c711101 (.i_clk(tick), .i_in(), .o_out(w711101));
	wire w171103;
	repeater #(1, 1'b1, 0, 0) c171103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171103));
	wire w331103;
	repeater #(1, 1'b0, 0, 0) c331103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w331103));
	wire w511103;
	repeater #(1, 1'b1, 0, 0) c511103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w511103));
	wire w671103;
	repeater #(1, 1'b0, 0, 0) c671103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w671103));
	wire w1811103;
	repeater #(1, 1'b0, 0, 0) c1811103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1811103));
	wire w301105;
	torch #(1'b1) c301105 (.i_clk(tick), .i_in(), .o_out(w301105));
	wire w641105;
	torch #(1'b1) c641105 (.i_clk(tick), .i_in(), .o_out(w641105));
	wire w1511105;
	repeater #(1, 1'b0, 0, 0) c1511105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1511105));
	wire w1841105;
	repeater #(1, 1'b1, 0, 0) c1841105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1841105));
	wire w221107;
	torch #(1'b1) c221107 (.i_clk(tick), .i_in(), .o_out(w221107));
	wire w381107;
	torch #(1'b1) c381107 (.i_clk(tick), .i_in(), .o_out(w381107));
	wire w561107;
	torch #(1'b1) c561107 (.i_clk(tick), .i_in(), .o_out(w561107));
	wire w721107;
	torch #(1'b1) c721107 (.i_clk(tick), .i_in(), .o_out(w721107));
	wire w291108;
	repeater #(1, 1'b0, 0, 0) c291108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w291108));
	wire w411108;
	repeater #(1, 1'b0, 0, 0) c411108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w411108));
	wire w631108;
	repeater #(1, 1'b0, 0, 0) c631108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w631108));
	wire w751108;
	repeater #(1, 1'b0, 0, 0) c751108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w751108));
	wire w1601108;
	torch #(1'b1) c1601108 (.i_clk(tick), .i_in(), .o_out(w1601108));
	wire w1641108;
	torch #(1'b1) c1641108 (.i_clk(tick), .i_in(), .o_out(w1641108));
	wire w1681108;
	torch #(1'b1) c1681108 (.i_clk(tick), .i_in(), .o_out(w1681108));
	wire w1721108;
	torch #(1'b1) c1721108 (.i_clk(tick), .i_in(), .o_out(w1721108));
	wire w231109;
	repeater #(1, 1'b0, 0, 0) c231109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w231109));
	wire w351109;
	repeater #(1, 1'b0, 0, 0) c351109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w351109));
	wire w571109;
	repeater #(1, 1'b0, 0, 0) c571109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w571109));
	wire w691109;
	repeater #(1, 1'b0, 0, 0) c691109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691109));
	wire w351111;
	repeater #(1, 1'b0, 0, 0) c351111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w351111));
	wire w691111;
	repeater #(1, 1'b0, 0, 0) c691111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691111));
	wire w1531112;
	torch #(1'b0) c1531112 (.i_clk(tick), .i_in(), .o_out(w1531112));
	wire w1571112;
	torch #(1'b0) c1571112 (.i_clk(tick), .i_in(), .o_out(w1571112));
	wire w1611112;
	torch #(1'b0) c1611112 (.i_clk(tick), .i_in(), .o_out(w1611112));
	wire w1651112;
	torch #(1'b1) c1651112 (.i_clk(tick), .i_in(), .o_out(w1651112));
	wire w1691112;
	torch #(1'b0) c1691112 (.i_clk(tick), .i_in(), .o_out(w1691112));
	wire w1731112;
	torch #(1'b0) c1731112 (.i_clk(tick), .i_in(), .o_out(w1731112));
	wire w1771112;
	torch #(1'b0) c1771112 (.i_clk(tick), .i_in(), .o_out(w1771112));
	wire w1541114;
	torch #(1'b1) c1541114 (.i_clk(tick), .i_in(), .o_out(w1541114));
	wire w1581114;
	torch #(1'b1) c1581114 (.i_clk(tick), .i_in(), .o_out(w1581114));
	wire w1621114;
	torch #(1'b1) c1621114 (.i_clk(tick), .i_in(), .o_out(w1621114));
	wire w1661114;
	torch #(1'b1) c1661114 (.i_clk(tick), .i_in(), .o_out(w1661114));
	wire w1701114;
	torch #(1'b1) c1701114 (.i_clk(tick), .i_in(), .o_out(w1701114));
	wire w1741114;
	torch #(1'b1) c1741114 (.i_clk(tick), .i_in(), .o_out(w1741114));
	wire w1781114;
	torch #(1'b1) c1781114 (.i_clk(tick), .i_in(), .o_out(w1781114));
	wire w1551116;
	torch #(1'b0) c1551116 (.i_clk(tick), .i_in(), .o_out(w1551116));
	wire w1591116;
	torch #(1'b0) c1591116 (.i_clk(tick), .i_in(), .o_out(w1591116));
	wire w1631116;
	torch #(1'b0) c1631116 (.i_clk(tick), .i_in(), .o_out(w1631116));
	wire w1671116;
	torch #(1'b0) c1671116 (.i_clk(tick), .i_in(), .o_out(w1671116));
	wire w1711116;
	torch #(1'b0) c1711116 (.i_clk(tick), .i_in(), .o_out(w1711116));
	wire w1751116;
	torch #(1'b0) c1751116 (.i_clk(tick), .i_in(), .o_out(w1751116));
	wire w1791116;
	torch #(1'b0) c1791116 (.i_clk(tick), .i_in(), .o_out(w1791116));
	wire w1811119;
	repeater #(1, 1'b0, 0, 0) c1811119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1811119));
	wire w1511121;
	repeater #(1, 1'b0, 0, 0) c1511121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1511121));
	wire w1841123;
	repeater #(1, 1'b1, 0, 0) c1841123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1841123));
	wire w1601124;
	torch #(1'b1) c1601124 (.i_clk(tick), .i_in(), .o_out(w1601124));
	wire w1641124;
	torch #(1'b1) c1641124 (.i_clk(tick), .i_in(), .o_out(w1641124));
	wire w1681124;
	torch #(1'b1) c1681124 (.i_clk(tick), .i_in(), .o_out(w1681124));
	wire w1721124;
	torch #(1'b1) c1721124 (.i_clk(tick), .i_in(), .o_out(w1721124));
	wire w1531128;
	torch #(1'b0) c1531128 (.i_clk(tick), .i_in(), .o_out(w1531128));
	wire w1571128;
	torch #(1'b0) c1571128 (.i_clk(tick), .i_in(), .o_out(w1571128));
	wire w1611128;
	torch #(1'b1) c1611128 (.i_clk(tick), .i_in(), .o_out(w1611128));
	wire w1651128;
	torch #(1'b0) c1651128 (.i_clk(tick), .i_in(), .o_out(w1651128));
	wire w1691128;
	torch #(1'b1) c1691128 (.i_clk(tick), .i_in(), .o_out(w1691128));
	wire w1731128;
	torch #(1'b0) c1731128 (.i_clk(tick), .i_in(), .o_out(w1731128));
	wire w1771128;
	torch #(1'b0) c1771128 (.i_clk(tick), .i_in(), .o_out(w1771128));
	wire w1541130;
	torch #(1'b1) c1541130 (.i_clk(tick), .i_in(), .o_out(w1541130));
	wire w1581130;
	torch #(1'b1) c1581130 (.i_clk(tick), .i_in(), .o_out(w1581130));
	wire w1621130;
	torch #(1'b1) c1621130 (.i_clk(tick), .i_in(), .o_out(w1621130));
	wire w1661130;
	torch #(1'b1) c1661130 (.i_clk(tick), .i_in(), .o_out(w1661130));
	wire w1701130;
	torch #(1'b1) c1701130 (.i_clk(tick), .i_in(), .o_out(w1701130));
	wire w1741130;
	torch #(1'b1) c1741130 (.i_clk(tick), .i_in(), .o_out(w1741130));
	wire w1781130;
	torch #(1'b1) c1781130 (.i_clk(tick), .i_in(), .o_out(w1781130));
	wire w1551132;
	torch #(1'b0) c1551132 (.i_clk(tick), .i_in(), .o_out(w1551132));
	wire w1591132;
	torch #(1'b0) c1591132 (.i_clk(tick), .i_in(), .o_out(w1591132));
	wire w1631132;
	torch #(1'b0) c1631132 (.i_clk(tick), .i_in(), .o_out(w1631132));
	wire w1671132;
	torch #(1'b0) c1671132 (.i_clk(tick), .i_in(), .o_out(w1671132));
	wire w1711132;
	torch #(1'b0) c1711132 (.i_clk(tick), .i_in(), .o_out(w1711132));
	wire w1751132;
	torch #(1'b0) c1751132 (.i_clk(tick), .i_in(), .o_out(w1751132));
	wire w1791132;
	torch #(1'b0) c1791132 (.i_clk(tick), .i_in(), .o_out(w1791132));
	wire w1811135;
	repeater #(1, 1'b0, 0, 0) c1811135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1811135));
	wire w13501;
	repeater #(1, 1'b0, 0, 0) c13501 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13501));
	wire w14404;
	torch #(1'b1) c14404 (.i_clk(tick), .i_in(), .o_out(w14404));
	wire w14804;
	torch #(1'b1) c14804 (.i_clk(tick), .i_in(), .o_out(w14804));
	wire w15204;
	torch #(1'b1) c15204 (.i_clk(tick), .i_in(), .o_out(w15204));
	wire w15604;
	torch #(1'b1) c15604 (.i_clk(tick), .i_in(), .o_out(w15604));
	wire w16805;
	repeater #(1, 1'b1, 0, 0) c16805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16805));
	wire w13708;
	torch #(1'b0) c13708 (.i_clk(tick), .i_in(), .o_out(w13708));
	wire w14108;
	torch #(1'b0) c14108 (.i_clk(tick), .i_in(), .o_out(w14108));
	wire w14508;
	torch #(1'b0) c14508 (.i_clk(tick), .i_in(), .o_out(w14508));
	wire w14908;
	torch #(1'b1) c14908 (.i_clk(tick), .i_in(), .o_out(w14908));
	wire w15308;
	torch #(1'b0) c15308 (.i_clk(tick), .i_in(), .o_out(w15308));
	wire w15708;
	torch #(1'b0) c15708 (.i_clk(tick), .i_in(), .o_out(w15708));
	wire w16108;
	torch #(1'b0) c16108 (.i_clk(tick), .i_in(), .o_out(w16108));
	wire w138010;
	torch #(1'b1) c138010 (.i_clk(tick), .i_in(), .o_out(w138010));
	wire w142010;
	torch #(1'b1) c142010 (.i_clk(tick), .i_in(), .o_out(w142010));
	wire w146010;
	torch #(1'b1) c146010 (.i_clk(tick), .i_in(), .o_out(w146010));
	wire w150010;
	torch #(1'b1) c150010 (.i_clk(tick), .i_in(), .o_out(w150010));
	wire w154010;
	torch #(1'b1) c154010 (.i_clk(tick), .i_in(), .o_out(w154010));
	wire w158010;
	torch #(1'b1) c158010 (.i_clk(tick), .i_in(), .o_out(w158010));
	wire w162010;
	torch #(1'b1) c162010 (.i_clk(tick), .i_in(), .o_out(w162010));
	wire w139012;
	torch #(1'b0) c139012 (.i_clk(tick), .i_in(), .o_out(w139012));
	wire w143012;
	torch #(1'b0) c143012 (.i_clk(tick), .i_in(), .o_out(w143012));
	wire w147012;
	torch #(1'b0) c147012 (.i_clk(tick), .i_in(), .o_out(w147012));
	wire w151012;
	torch #(1'b0) c151012 (.i_clk(tick), .i_in(), .o_out(w151012));
	wire w155012;
	torch #(1'b0) c155012 (.i_clk(tick), .i_in(), .o_out(w155012));
	wire w159012;
	torch #(1'b0) c159012 (.i_clk(tick), .i_in(), .o_out(w159012));
	wire w163012;
	torch #(1'b0) c163012 (.i_clk(tick), .i_in(), .o_out(w163012));
	wire w169020;

	wire w170020;

	wire w168022;
	repeater #(1, 1'b1, 0, 0) c168022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168022));
	wire w171022;
	repeater #(1, 1'b0, 0, 0) c171022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171022));
	wire w148023;
	repeater #(1, 1'b1, 0, 0) c148023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148023));
	wire w165024;
	repeater #(1, 1'b1, 0, 0) c165024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165024));
	wire w149027;
	repeater #(1, 1'b1, 0, 0) c149027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149027));
	wire w161027;
	repeater #(1, 1'b1, 0, 0) c161027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161027));
	wire w171028;
	torch #(1'b1) c171028 (.i_clk(tick), .i_in(), .o_out(w171028));
	wire w169029;
	torch #(1'b0) c169029 (.i_clk(tick), .i_in(), .o_out(w169029));
	wire w26071;

	wire w59071;

	wire w60071;

	wire w93071;

	wire w94071;

	wire w127071;

	wire w128071;

	wire w161071;

	wire w27072;
	repeater #(1, 1'b1, 0, 0) c27072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27072));
	wire w61072;
	repeater #(1, 1'b1, 0, 0) c61072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61072));
	wire w95072;
	repeater #(1, 1'b1, 0, 0) c95072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95072));
	wire w129072;
	repeater #(1, 1'b1, 0, 0) c129072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w129072));
	wire w24073;

	wire w57073;

	wire w58073;

	wire w91073;

	wire w92073;

	wire w125073;

	wire w126073;

	wire w159073;

	wire w162073;
	repeater #(1, 1'b1, 0, 0) c162073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162073));
	wire w25074;
	repeater #(1, 1'b1, 0, 0) c25074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25074));
	wire w59074;
	repeater #(1, 1'b1, 0, 0) c59074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59074));
	wire w93074;
	repeater #(1, 1'b1, 0, 0) c93074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93074));
	wire w127074;
	repeater #(1, 1'b1, 0, 0) c127074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127074));
	wire w161074;

	wire w22075;

	wire w55075;

	wire w56075;

	wire w89075;

	wire w90075;

	wire w123075;

	wire w124075;

	wire w157075;

	wire w160075;
	repeater #(1, 1'b1, 0, 0) c160075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160075));
	wire w23076;
	repeater #(1, 1'b1, 0, 0) c23076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23076));
	wire w57076;
	repeater #(1, 1'b1, 0, 0) c57076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57076));
	wire w91076;
	repeater #(1, 1'b1, 0, 0) c91076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91076));
	wire w125076;
	repeater #(1, 1'b1, 0, 0) c125076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125076));
	wire w159076;

	wire w20077;

	wire w53077;

	wire w54077;

	wire w87077;

	wire w88077;

	wire w121077;

	wire w122077;

	wire w155077;

	wire w158077;
	repeater #(1, 1'b1, 0, 0) c158077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158077));
	wire w21078;
	repeater #(1, 1'b1, 0, 0) c21078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21078));
	wire w55078;
	repeater #(1, 1'b1, 0, 0) c55078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55078));
	wire w89078;
	repeater #(1, 1'b1, 0, 0) c89078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89078));
	wire w123078;
	repeater #(1, 1'b1, 0, 0) c123078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123078));
	wire w157078;

	wire w18079;

	wire w51079;

	wire w52079;

	wire w85079;

	wire w86079;

	wire w119079;

	wire w120079;

	wire w153079;

	wire w156079;
	repeater #(1, 1'b1, 0, 0) c156079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156079));
	wire w19080;
	repeater #(1, 1'b0, 0, 0) c19080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19080));
	wire w53080;
	repeater #(1, 1'b0, 0, 0) c53080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53080));
	wire w87080;
	repeater #(1, 1'b0, 0, 0) c87080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87080));
	wire w121080;
	repeater #(1, 1'b0, 0, 0) c121080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121080));
	wire w155080;

	wire w16081;

	wire w49081;

	wire w50081;

	wire w83081;

	wire w84081;

	wire w117081;

	wire w118081;

	wire w151081;

	wire w154081;
	repeater #(1, 1'b0, 0, 0) c154081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154081));
	wire w17082;
	repeater #(1, 1'b0, 0, 0) c17082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17082));
	wire w51082;
	repeater #(1, 1'b0, 0, 0) c51082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51082));
	wire w85082;
	repeater #(1, 1'b0, 0, 0) c85082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85082));
	wire w119082;
	repeater #(1, 1'b0, 0, 0) c119082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119082));
	wire w153082;

	wire w14083;

	wire w47083;

	wire w48083;

	wire w81083;

	wire w82083;

	wire w115083;

	wire w116083;

	wire w149083;

	wire w152083;
	repeater #(1, 1'b0, 0, 0) c152083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152083));
	wire w15084;
	repeater #(1, 1'b1, 0, 0) c15084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15084));
	wire w49084;
	repeater #(1, 1'b1, 0, 0) c49084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49084));
	wire w83084;
	repeater #(1, 1'b1, 0, 0) c83084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83084));
	wire w117084;
	repeater #(1, 1'b1, 0, 0) c117084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117084));
	wire w151084;

	wire w12085;

	wire w45085;

	wire w46085;

	wire w79085;

	wire w80085;

	wire w113085;

	wire w114085;

	wire w147085;

	wire w150085;
	repeater #(1, 1'b1, 0, 0) c150085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150085));
	wire w13086;
	repeater #(1, 1'b0, 0, 0) c13086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13086));
	wire w47086;
	repeater #(1, 1'b0, 0, 0) c47086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47086));
	wire w81086;
	repeater #(1, 1'b0, 0, 0) c81086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81086));
	wire w115086;
	repeater #(1, 1'b0, 0, 0) c115086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115086));
	wire w149086;

	wire w10087;

	wire w43087;

	wire w44087;

	wire w77087;

	wire w78087;

	wire w111087;

	wire w112087;

	wire w145087;

	wire w148087;
	repeater #(1, 1'b0, 0, 0) c148087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148087));
	wire w11088;
	repeater #(1, 1'b0, 0, 0) c11088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11088));
	wire w45088;
	repeater #(1, 1'b0, 0, 0) c45088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45088));
	wire w79088;
	repeater #(1, 1'b0, 0, 0) c79088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79088));
	wire w113088;
	repeater #(1, 1'b0, 0, 0) c113088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113088));
	wire w147088;

	wire w8089;

	wire w41089;

	wire w42089;

	wire w75089;

	wire w76089;

	wire w109089;

	wire w110089;

	wire w143089;

	wire w146089;
	repeater #(1, 1'b0, 0, 0) c146089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146089));
	wire w9090;
	repeater #(1, 1'b0, 0, 0) c9090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9090));
	wire w43090;
	repeater #(1, 1'b0, 0, 0) c43090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43090));
	wire w77090;
	repeater #(1, 1'b0, 0, 0) c77090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77090));
	wire w111090;
	repeater #(1, 1'b0, 0, 0) c111090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111090));
	wire w145090;

	wire w6091;

	wire w39091;

	wire w40091;

	wire w73091;

	wire w74091;

	wire w107091;

	wire w108091;

	wire w141091;

	wire w144091;
	repeater #(1, 1'b0, 0, 0) c144091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144091));
	wire w7092;
	repeater #(1, 1'b1, 0, 0) c7092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7092));
	wire w41092;
	repeater #(1, 1'b1, 0, 0) c41092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41092));
	wire w75092;
	repeater #(1, 1'b1, 0, 0) c75092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75092));
	wire w109092;
	repeater #(1, 1'b1, 0, 0) c109092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109092));
	wire w143092;

	wire w4093;

	wire w37093;

	wire w38093;

	wire w71093;

	wire w72093;

	wire w105093;

	wire w106093;

	wire w139093;

	wire w142093;
	repeater #(1, 1'b1, 0, 0) c142093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142093));
	wire w5094;
	repeater #(1, 1'b1, 0, 0) c5094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5094));
	wire w39094;
	repeater #(1, 1'b1, 0, 0) c39094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39094));
	wire w73094;
	repeater #(1, 1'b1, 0, 0) c73094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73094));
	wire w107094;
	repeater #(1, 1'b1, 0, 0) c107094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107094));
	wire w141094;

	wire w2095;

	wire w35095;

	wire w36095;

	wire w69095;

	wire w70095;

	wire w103095;

	wire w104095;

	wire w137095;

	wire w140095;
	repeater #(1, 1'b1, 0, 0) c140095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140095));
	wire w3096;
	repeater #(1, 1'b1, 0, 0) c3096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3096));
	wire w37096;
	repeater #(1, 1'b1, 0, 0) c37096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37096));
	wire w71096;
	repeater #(1, 1'b1, 0, 0) c71096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71096));
	wire w105096;
	repeater #(1, 1'b1, 0, 0) c105096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105096));
	wire w139096;

	wire w33097;

	wire w67097;

	wire w101097;

	wire w135097;

	wire w138097;
	repeater #(1, 1'b1, 0, 0) c138097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138097));
	wire w1098;
	repeater #(1, 1'b1, 0, 0) c1098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1098));
	wire w35098;
	repeater #(1, 1'b1, 0, 0) c35098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35098));
	wire w69098;
	repeater #(1, 1'b1, 0, 0) c69098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69098));
	wire w103098;
	repeater #(1, 1'b1, 0, 0) c103098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103098));
	wire w137098;

	wire w136099;
	repeater #(2, 1'b1, 0, 0) c136099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136099));
	wire w1380100;
	repeater #(1, 1'b1, 0, 0) c1380100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380100));
	wire w200103;
	repeater #(2, 1'b1, 0, 0) c200103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200103));
	wire w540103;
	repeater #(2, 1'b1, 0, 0) c540103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540103));
	wire w1370103;
	torch #(1'b1) c1370103 (.i_clk(tick), .i_in(), .o_out(w1370103));
	wire w1410103;
	torch #(1'b1) c1410103 (.i_clk(tick), .i_in(), .o_out(w1410103));
	wire w1450103;
	torch #(1'b1) c1450103 (.i_clk(tick), .i_in(), .o_out(w1450103));
	wire w1490103;
	torch #(1'b0) c1490103 (.i_clk(tick), .i_in(), .o_out(w1490103));
	wire w1530103;
	torch #(1'b1) c1530103 (.i_clk(tick), .i_in(), .o_out(w1530103));
	wire w1570103;
	torch #(1'b1) c1570103 (.i_clk(tick), .i_in(), .o_out(w1570103));
	wire w1610103;
	torch #(1'b1) c1610103 (.i_clk(tick), .i_in(), .o_out(w1610103));
	wire w60105;
	repeater #(1, 1'b1, 0, 0) c60105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60105));
	wire w120105;
	torch #(1'b0) c120105 (.i_clk(tick), .i_in(), .o_out(w120105));
	wire w220105;
	repeater #(1, 1'b1, 0, 0) c220105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220105));
	wire w400105;
	repeater #(1, 1'b1, 0, 0) c400105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400105));
	wire w460105;
	torch #(1'b0) c460105 (.i_clk(tick), .i_in(), .o_out(w460105));
	wire w560105;
	repeater #(1, 1'b1, 0, 0) c560105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560105));
	wire w1380106;
	repeater #(1, 1'b1, 0, 0) c1380106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380106));
	wire w1420106;
	repeater #(1, 1'b1, 0, 0) c1420106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420106));
	wire w1460106;
	repeater #(1, 1'b1, 0, 0) c1460106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460106));
	wire w1500106;
	repeater #(1, 1'b0, 0, 0) c1500106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500106));
	wire w1540106;
	repeater #(1, 1'b1, 0, 0) c1540106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540106));
	wire w1580106;
	repeater #(1, 1'b1, 0, 0) c1580106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580106));
	wire w1620106;
	repeater #(1, 1'b1, 0, 0) c1620106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620106));
	wire w1370107;
	torch #(1'b1) c1370107 (.i_clk(tick), .i_in(), .o_out(w1370107));
	wire w1410107;
	torch #(1'b1) c1410107 (.i_clk(tick), .i_in(), .o_out(w1410107));
	wire w1450107;
	torch #(1'b1) c1450107 (.i_clk(tick), .i_in(), .o_out(w1450107));
	wire w1490107;
	torch #(1'b0) c1490107 (.i_clk(tick), .i_in(), .o_out(w1490107));
	wire w1530107;
	torch #(1'b1) c1530107 (.i_clk(tick), .i_in(), .o_out(w1530107));
	wire w1570107;
	torch #(1'b1) c1570107 (.i_clk(tick), .i_in(), .o_out(w1570107));
	wire w1610107;
	torch #(1'b1) c1610107 (.i_clk(tick), .i_in(), .o_out(w1610107));
	wire w130108;
	repeater #(1, 1'b1, 0, 0) c130108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130108));
	wire w470108;
	repeater #(1, 1'b0, 0, 0) c470108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470108));
	wire w60109;
	repeater #(1, 1'b1, 0, 0) c60109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60109));
	wire w220109;
	repeater #(1, 1'b1, 0, 0) c220109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220109));
	wire w400109;
	repeater #(1, 1'b1, 0, 0) c400109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400109));
	wire w560109;
	repeater #(1, 1'b1, 0, 0) c560109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560109));
	wire w110110;

	wire w450110;

	wire w1360110;
	torch #(1'b0) c1360110 (.i_clk(tick), .i_in(), .o_out(w1360110));
	wire w1400110;
	torch #(1'b0) c1400110 (.i_clk(tick), .i_in(), .o_out(w1400110));
	wire w1440110;
	torch #(1'b1) c1440110 (.i_clk(tick), .i_in(), .o_out(w1440110));
	wire w1480110;
	torch #(1'b1) c1480110 (.i_clk(tick), .i_in(), .o_out(w1480110));
	wire w1520110;
	torch #(1'b1) c1520110 (.i_clk(tick), .i_in(), .o_out(w1520110));
	wire w1560110;
	torch #(1'b0) c1560110 (.i_clk(tick), .i_in(), .o_out(w1560110));
	wire w1600110;
	torch #(1'b0) c1600110 (.i_clk(tick), .i_in(), .o_out(w1600110));
	wire w30111;

	wire w190111;

	wire w370111;

	wire w530111;

	wire w00112;

	wire w50112;

	wire w60112;

	wire w160112;

	wire w220112;

	wire w340112;

	wire w390112;

	wire w400112;

	wire w500112;

	wire w560112;

	wire w2060113;

	wire w140114;

	wire w320114;

	wire w480114;

	wire w40115;

	wire w50115;

	wire w200115;

	wire w210115;

	wire w380115;

	wire w390115;

	wire w540115;

	wire w550115;

	wire w140116;

	wire w480116;

	wire w2060117;

	wire w20118;

	wire w60118;

	wire w100118;

	wire w140118;

	wire w180118;

	wire w220118;

	wire w320118;

	wire w360118;

	wire w400118;

	wire w440118;

	wire w480118;

	wire w520118;

	wire w560118;

	wire w2060121;

	wire w20122;

	wire w60122;

	wire w100122;

	wire w140122;

	wire w180122;

	wire w220122;

	wire w320122;

	wire w360122;

	wire w400122;

	wire w440122;

	wire w480122;

	wire w520122;

	wire w560122;

	wire w2040123;
	repeater #(1, 1'b1, 0, 0) c2040123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040123));
	wire w00124;
	repeater #(1, 1'b1, 0, 0) c00124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w00124));
	wire w40124;
	repeater #(1, 1'b1, 0, 0) c40124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40124));
	wire w80124;
	repeater #(1, 1'b1, 0, 0) c80124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80124));
	wire w300124;
	repeater #(1, 1'b1, 0, 0) c300124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300124));
	wire w340124;
	repeater #(1, 1'b1, 0, 0) c340124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340124));
	wire w380124;
	repeater #(1, 1'b1, 0, 0) c380124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380124));
	wire w420124;
	repeater #(1, 1'b0, 0, 0) c420124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420124));
	wire w140125;

	wire w180125;

	wire w220125;

	wire w480125;

	wire w520125;

	wire w560125;

	wire w1370125;
	torch #(1'b1) c1370125 (.i_clk(tick), .i_in(), .o_out(w1370125));
	wire w1410125;
	torch #(1'b1) c1410125 (.i_clk(tick), .i_in(), .o_out(w1410125));
	wire w1450125;
	torch #(1'b1) c1450125 (.i_clk(tick), .i_in(), .o_out(w1450125));
	wire w1490125;
	torch #(1'b0) c1490125 (.i_clk(tick), .i_in(), .o_out(w1490125));
	wire w1530125;
	torch #(1'b1) c1530125 (.i_clk(tick), .i_in(), .o_out(w1530125));
	wire w1570125;
	torch #(1'b1) c1570125 (.i_clk(tick), .i_in(), .o_out(w1570125));
	wire w1610125;
	torch #(1'b1) c1610125 (.i_clk(tick), .i_in(), .o_out(w1610125));
	wire w1380126;
	repeater #(1, 1'b0, 0, 0) c1380126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380126));
	wire w1420126;
	repeater #(1, 1'b0, 0, 0) c1420126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420126));
	wire w1460126;
	repeater #(1, 1'b1, 0, 0) c1460126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460126));
	wire w1500126;
	repeater #(1, 1'b1, 0, 0) c1500126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500126));
	wire w1540126;
	repeater #(1, 1'b1, 0, 0) c1540126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540126));
	wire w1580126;
	repeater #(1, 1'b0, 0, 0) c1580126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580126));
	wire w1620126;
	repeater #(1, 1'b0, 0, 0) c1620126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620126));
	wire w140127;

	wire w480127;

	wire w120128;
	repeater #(1, 1'b1, 0, 0) c120128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120128));
	wire w460128;
	repeater #(1, 1'b1, 0, 0) c460128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460128));
	wire w1360128;

	wire w1380128;
	repeater #(1, 1'b0, 0, 0) c1380128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380128));
	wire w1400128;

	wire w1420128;
	repeater #(1, 1'b0, 0, 0) c1420128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420128));
	wire w1440128;

	wire w1460128;
	repeater #(1, 1'b1, 0, 0) c1460128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460128));
	wire w1480128;

	wire w1500128;
	repeater #(1, 1'b1, 0, 0) c1500128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500128));
	wire w1520128;

	wire w1540128;
	repeater #(1, 1'b1, 0, 0) c1540128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540128));
	wire w1560128;

	wire w1580128;
	repeater #(1, 1'b0, 0, 0) c1580128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580128));
	wire w1600128;

	wire w1620128;
	repeater #(1, 1'b0, 0, 0) c1620128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620128));
	wire w30129;
	repeater #(1, 1'b1, 0, 0) c30129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30129));
	wire w190129;
	repeater #(1, 1'b1, 0, 0) c190129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190129));
	wire w370129;
	repeater #(1, 1'b1, 0, 0) c370129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370129));
	wire w530129;
	repeater #(1, 1'b1, 0, 0) c530129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530129));
	wire w2060129;

	wire w140130;

	wire w320130;

	wire w480130;

	wire w60131;

	wire w400131;

	wire w10132;

	wire w30132;

	wire w40132;

	wire w90132;

	wire w170132;

	wire w190132;

	wire w200132;

	wire w350132;

	wire w370132;

	wire w380132;

	wire w430132;

	wire w510132;

	wire w530132;

	wire w540132;

	wire w110134;

	wire w120134;

	wire w450134;

	wire w460134;

	wire w10136;

	wire w30136;

	wire w40136;

	wire w170136;

	wire w190136;

	wire w200136;

	wire w350136;

	wire w370136;

	wire w380136;

	wire w510136;

	wire w530136;

	wire w540136;

	wire w700137;
	repeater #(2, 1'b0, 0, 0) c700137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w700137));
	wire w750137;
	repeater #(2, 1'b0, 0, 0) c750137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w750137));
	wire w1230137;
	repeater #(2, 1'b0, 0, 0) c1230137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230137));
	wire w1280137;
	repeater #(2, 1'b0, 0, 0) c1280137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1280137));
	wire w2060137;
	torch #(1'b1) c2060137 (.i_clk(tick), .i_in(), .o_out(w2060137));
	wire w2070137;

	wire w140138;
	torch #(1'b1) c140138 (.i_clk(tick), .i_in(), .o_out(w140138));
	wire w150138;

	wire w200138;

	wire w320138;
	torch #(1'b1) c320138 (.i_clk(tick), .i_in(), .o_out(w320138));
	wire w330138;

	wire w480138;
	torch #(1'b1) c480138 (.i_clk(tick), .i_in(), .o_out(w480138));
	wire w490138;

	wire w540138;

	wire w2070138;

	wire w10139;

	wire w150139;

	wire w170139;

	wire w330139;

	wire w350139;

	wire w490139;

	wire w510139;

	wire w700139;

	wire w710139;

	wire w1270139;

	wire w1280139;

	wire w740140;
	repeater #(2, 1'b0, 0, 0) c740140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w740140));
	wire w750140;
	repeater #(2, 1'b0, 0, 0) c750140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w750140));
	wire w770140;

	wire w1210140;

	wire w1230140;
	repeater #(2, 1'b0, 0, 0) c1230140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230140));
	wire w1240140;
	repeater #(2, 1'b0, 0, 0) c1240140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240140));
	wire w10141;

	wire w20141;

	wire w30141;

	wire w170141;

	wire w180141;

	wire w190141;

	wire w350141;

	wire w360141;

	wire w370141;

	wire w510141;

	wire w520141;

	wire w530141;

	wire w750141;

	wire w770141;
	repeater #(1, 1'b0, 0, 0) c770141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w770141));
	wire w1210141;
	repeater #(1, 1'b0, 0, 0) c1210141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1210141));
	wire w1230141;

	wire w1370141;
	torch #(1'b1) c1370141 (.i_clk(tick), .i_in(), .o_out(w1370141));
	wire w1410141;
	torch #(1'b1) c1410141 (.i_clk(tick), .i_in(), .o_out(w1410141));
	wire w1450141;
	torch #(1'b0) c1450141 (.i_clk(tick), .i_in(), .o_out(w1450141));
	wire w1490141;
	torch #(1'b1) c1490141 (.i_clk(tick), .i_in(), .o_out(w1490141));
	wire w1530141;
	torch #(1'b0) c1530141 (.i_clk(tick), .i_in(), .o_out(w1530141));
	wire w1570141;
	torch #(1'b1) c1570141 (.i_clk(tick), .i_in(), .o_out(w1570141));
	wire w1610141;
	torch #(1'b1) c1610141 (.i_clk(tick), .i_in(), .o_out(w1610141));
	wire w30142;

	wire w120142;

	wire w130142;

	wire w190142;

	wire w370142;

	wire w460142;

	wire w470142;

	wire w530142;

	wire w710142;

	wire w750142;

	wire w1230142;

	wire w1270142;

	wire w1380142;
	repeater #(1, 1'b0, 0, 0) c1380142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380142));
	wire w1420142;
	repeater #(1, 1'b0, 0, 0) c1420142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420142));
	wire w1460142;
	repeater #(1, 1'b1, 0, 0) c1460142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460142));
	wire w1500142;
	repeater #(1, 1'b1, 0, 0) c1500142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500142));
	wire w1540142;
	repeater #(1, 1'b1, 0, 0) c1540142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540142));
	wire w1580142;
	repeater #(1, 1'b0, 0, 0) c1580142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580142));
	wire w1620142;
	repeater #(1, 1'b0, 0, 0) c1620142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620142));
	wire w710143;

	wire w730143;
	repeater #(1, 1'b0, 0, 0) c730143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w730143));
	wire w780143;

	wire w820143;

	wire w1160143;

	wire w1200143;

	wire w1250143;
	repeater #(1, 1'b0, 0, 0) c1250143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1250143));
	wire w1270143;

	wire w10144;
	repeater #(1, 1'b0, 0, 0) c10144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10144));
	wire w30144;
	torch #(1'b0) c30144 (.i_clk(tick), .i_in(), .o_out(w30144));
	wire w90144;
	torch #(1'b0) c90144 (.i_clk(tick), .i_in(), .o_out(w90144));
	wire w170144;
	repeater #(1, 1'b0, 0, 0) c170144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170144));
	wire w190144;
	torch #(1'b0) c190144 (.i_clk(tick), .i_in(), .o_out(w190144));
	wire w250144;
	torch #(1'b0) c250144 (.i_clk(tick), .i_in(), .o_out(w250144));
	wire w350144;
	repeater #(1, 1'b0, 0, 0) c350144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w350144));
	wire w370144;
	torch #(1'b0) c370144 (.i_clk(tick), .i_in(), .o_out(w370144));
	wire w430144;
	torch #(1'b0) c430144 (.i_clk(tick), .i_in(), .o_out(w430144));
	wire w510144;
	repeater #(1, 1'b0, 0, 0) c510144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510144));
	wire w530144;
	torch #(1'b0) c530144 (.i_clk(tick), .i_in(), .o_out(w530144));
	wire w590144;
	torch #(1'b0) c590144 (.i_clk(tick), .i_in(), .o_out(w590144));
	wire w780144;

	wire w800144;
	repeater #(1, 1'b0, 0, 0) c800144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800144));
	wire w810144;

	wire w1170144;

	wire w1180144;
	repeater #(1, 1'b0, 0, 0) c1180144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1180144));
	wire w1200144;

	wire w1360144;

	wire w1380144;
	repeater #(1, 1'b0, 0, 0) c1380144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380144));
	wire w1400144;

	wire w1420144;
	repeater #(1, 1'b0, 0, 0) c1420144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420144));
	wire w1440144;

	wire w1460144;
	repeater #(1, 1'b1, 0, 0) c1460144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460144));
	wire w1480144;

	wire w1500144;
	repeater #(1, 1'b1, 0, 0) c1500144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500144));
	wire w1520144;

	wire w1540144;
	repeater #(1, 1'b1, 0, 0) c1540144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540144));
	wire w1560144;

	wire w1580144;
	repeater #(1, 1'b0, 0, 0) c1580144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580144));
	wire w1600144;

	wire w1620144;
	repeater #(1, 1'b0, 0, 0) c1620144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620144));
	wire w740145;

	wire w1240145;

	wire w50146;
	repeater #(1, 1'b1, 0, 0) c50146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50146));
	wire w210146;
	repeater #(1, 1'b1, 0, 0) c210146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210146));
	wire w390146;
	repeater #(1, 1'b1, 0, 0) c390146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390146));
	wire w550146;
	repeater #(1, 1'b1, 0, 0) c550146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550146));
	wire w710146;

	wire w720146;
	repeater #(1, 1'b0, 0, 0) c720146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w720146));
	wire w790146;
	repeater #(2, 1'b0, 0, 0) c790146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w790146));
	wire w1190146;
	repeater #(2, 1'b0, 0, 0) c1190146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190146));
	wire w1260146;
	repeater #(1, 1'b0, 0, 0) c1260146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1260146));
	wire w1270146;

	wire w20148;
	torch #(1'b1) c20148 (.i_clk(tick), .i_in(), .o_out(w20148));
	wire w180148;
	torch #(1'b1) c180148 (.i_clk(tick), .i_in(), .o_out(w180148));
	wire w360148;
	torch #(1'b1) c360148 (.i_clk(tick), .i_in(), .o_out(w360148));
	wire w520148;
	torch #(1'b1) c520148 (.i_clk(tick), .i_in(), .o_out(w520148));
	wire w100150;
	torch #(1'b1) c100150 (.i_clk(tick), .i_in(), .o_out(w100150));
	wire w260150;
	torch #(1'b1) c260150 (.i_clk(tick), .i_in(), .o_out(w260150));
	wire w440150;
	torch #(1'b1) c440150 (.i_clk(tick), .i_in(), .o_out(w440150));
	wire w600150;
	torch #(1'b1) c600150 (.i_clk(tick), .i_in(), .o_out(w600150));
	wire w10151;
	repeater #(1, 1'b0, 0, 0) c10151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10151));
	wire w170151;
	repeater #(1, 1'b0, 0, 0) c170151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170151));
	wire w350151;
	repeater #(1, 1'b0, 0, 0) c350151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w350151));
	wire w510151;
	repeater #(1, 1'b0, 0, 0) c510151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510151));
	wire w110152;
	repeater #(1, 1'b0, 0, 0) c110152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110152));
	wire w230152;
	repeater #(1, 1'b0, 0, 0) c230152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230152));
	wire w450152;
	repeater #(1, 1'b0, 0, 0) c450152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w450152));
	wire w570152;
	repeater #(1, 1'b0, 0, 0) c570152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570152));
	wire w230154;
	repeater #(1, 1'b0, 0, 0) c230154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230154));
	wire w570154;
	repeater #(1, 1'b0, 0, 0) c570154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570154));
	wire w1370157;
	torch #(1'b1) c1370157 (.i_clk(tick), .i_in(), .o_out(w1370157));
	wire w1410157;
	torch #(1'b1) c1410157 (.i_clk(tick), .i_in(), .o_out(w1410157));
	wire w1450157;
	torch #(1'b1) c1450157 (.i_clk(tick), .i_in(), .o_out(w1450157));
	wire w1490157;
	torch #(1'b0) c1490157 (.i_clk(tick), .i_in(), .o_out(w1490157));
	wire w1530157;
	torch #(1'b1) c1530157 (.i_clk(tick), .i_in(), .o_out(w1530157));
	wire w1570157;
	torch #(1'b1) c1570157 (.i_clk(tick), .i_in(), .o_out(w1570157));
	wire w1610157;
	torch #(1'b1) c1610157 (.i_clk(tick), .i_in(), .o_out(w1610157));
	wire w1380158;
	repeater #(1, 1'b0, 0, 0) c1380158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380158));
	wire w1420158;
	repeater #(1, 1'b0, 0, 0) c1420158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420158));
	wire w1460158;
	repeater #(1, 1'b1, 0, 0) c1460158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460158));
	wire w1500158;
	repeater #(1, 1'b1, 0, 0) c1500158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500158));
	wire w1540158;
	repeater #(1, 1'b1, 0, 0) c1540158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540158));
	wire w1580158;
	repeater #(1, 1'b0, 0, 0) c1580158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580158));
	wire w1620158;
	repeater #(1, 1'b0, 0, 0) c1620158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620158));
	wire w1360160;

	wire w1380160;
	repeater #(1, 1'b0, 0, 0) c1380160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380160));
	wire w1400160;

	wire w1420160;
	repeater #(1, 1'b0, 0, 0) c1420160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420160));
	wire w1440160;

	wire w1460160;
	repeater #(1, 1'b1, 0, 0) c1460160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460160));
	wire w1480160;

	wire w1500160;
	repeater #(1, 1'b1, 0, 0) c1500160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500160));
	wire w1520160;

	wire w1540160;
	repeater #(1, 1'b1, 0, 0) c1540160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540160));
	wire w1560160;

	wire w1580160;
	repeater #(1, 1'b0, 0, 0) c1580160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580160));
	wire w1600160;

	wire w1620160;
	repeater #(1, 1'b0, 0, 0) c1620160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620160));
	wire w1370173;
	torch #(1'b1) c1370173 (.i_clk(tick), .i_in(), .o_out(w1370173));
	wire w1410173;
	torch #(1'b1) c1410173 (.i_clk(tick), .i_in(), .o_out(w1410173));
	wire w1450173;
	torch #(1'b0) c1450173 (.i_clk(tick), .i_in(), .o_out(w1450173));
	wire w1490173;
	torch #(1'b1) c1490173 (.i_clk(tick), .i_in(), .o_out(w1490173));
	wire w1530173;
	torch #(1'b0) c1530173 (.i_clk(tick), .i_in(), .o_out(w1530173));
	wire w1570173;
	torch #(1'b1) c1570173 (.i_clk(tick), .i_in(), .o_out(w1570173));
	wire w1610173;
	torch #(1'b1) c1610173 (.i_clk(tick), .i_in(), .o_out(w1610173));
	wire w1380174;
	repeater #(1, 1'b0, 0, 0) c1380174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380174));
	wire w1420174;
	repeater #(1, 1'b0, 0, 0) c1420174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420174));
	wire w1460174;
	repeater #(1, 1'b1, 0, 0) c1460174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460174));
	wire w1500174;
	repeater #(1, 1'b1, 0, 0) c1500174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500174));
	wire w1540174;
	repeater #(1, 1'b1, 0, 0) c1540174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540174));
	wire w1580174;
	repeater #(1, 1'b0, 0, 0) c1580174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580174));
	wire w1620174;
	repeater #(1, 1'b0, 0, 0) c1620174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620174));
	wire w1360176;

	wire w1380176;
	repeater #(1, 1'b0, 0, 0) c1380176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380176));
	wire w1400176;

	wire w1420176;
	repeater #(1, 1'b0, 0, 0) c1420176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420176));
	wire w1440176;

	wire w1460176;
	repeater #(1, 1'b1, 0, 0) c1460176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460176));
	wire w1480176;

	wire w1500176;
	repeater #(1, 1'b1, 0, 0) c1500176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500176));
	wire w1520176;

	wire w1540176;
	repeater #(1, 1'b1, 0, 0) c1540176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540176));
	wire w1560176;

	wire w1580176;
	repeater #(1, 1'b0, 0, 0) c1580176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580176));
	wire w1600176;

	wire w1620176;
	repeater #(1, 1'b0, 0, 0) c1620176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620176));
	wire w137110;
	torch #(1'b1) c137110 (.i_clk(tick), .i_in(), .o_out(w137110));
	wire w141110;
	torch #(1'b1) c141110 (.i_clk(tick), .i_in(), .o_out(w141110));
	wire w145110;
	torch #(1'b1) c145110 (.i_clk(tick), .i_in(), .o_out(w145110));
	wire w149110;
	torch #(1'b0) c149110 (.i_clk(tick), .i_in(), .o_out(w149110));
	wire w153110;
	torch #(1'b1) c153110 (.i_clk(tick), .i_in(), .o_out(w153110));
	wire w157110;
	torch #(1'b1) c157110 (.i_clk(tick), .i_in(), .o_out(w157110));
	wire w161110;
	torch #(1'b1) c161110 (.i_clk(tick), .i_in(), .o_out(w161110));
	wire w138111;
	repeater #(1, 1'b0, 0, 0) c138111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138111));
	wire w142111;
	repeater #(1, 1'b0, 0, 0) c142111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142111));
	wire w146111;
	repeater #(1, 1'b1, 0, 0) c146111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146111));
	wire w150111;
	repeater #(1, 1'b1, 0, 0) c150111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150111));
	wire w154111;
	repeater #(1, 1'b1, 0, 0) c154111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154111));
	wire w158111;
	repeater #(1, 1'b0, 0, 0) c158111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158111));
	wire w162111;
	repeater #(1, 1'b0, 0, 0) c162111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162111));
	wire w136113;

	wire w138113;
	repeater #(1, 1'b0, 0, 0) c138113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138113));
	wire w140113;

	wire w142113;
	repeater #(1, 1'b0, 0, 0) c142113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142113));
	wire w144113;

	wire w146113;
	repeater #(1, 1'b1, 0, 0) c146113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146113));
	wire w148113;

	wire w150113;
	repeater #(1, 1'b1, 0, 0) c150113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150113));
	wire w152113;

	wire w154113;
	repeater #(1, 1'b1, 0, 0) c154113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154113));
	wire w156113;

	wire w158113;
	repeater #(1, 1'b0, 0, 0) c158113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158113));
	wire w160113;

	wire w162113;
	repeater #(1, 1'b0, 0, 0) c162113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162113));
	wire w137119;
	torch #(1'b1) c137119 (.i_clk(tick), .i_in(), .o_out(w137119));
	wire w141119;
	torch #(1'b1) c141119 (.i_clk(tick), .i_in(), .o_out(w141119));
	wire w145119;
	torch #(1'b0) c145119 (.i_clk(tick), .i_in(), .o_out(w145119));
	wire w149119;
	torch #(1'b0) c149119 (.i_clk(tick), .i_in(), .o_out(w149119));
	wire w153119;
	torch #(1'b0) c153119 (.i_clk(tick), .i_in(), .o_out(w153119));
	wire w157119;
	torch #(1'b1) c157119 (.i_clk(tick), .i_in(), .o_out(w157119));
	wire w161119;
	torch #(1'b1) c161119 (.i_clk(tick), .i_in(), .o_out(w161119));
	wire w136128;
	torch #(1'b1) c136128 (.i_clk(tick), .i_in(), .o_out(w136128));
	wire w140128;
	torch #(1'b1) c140128 (.i_clk(tick), .i_in(), .o_out(w140128));
	wire w144128;
	torch #(1'b1) c144128 (.i_clk(tick), .i_in(), .o_out(w144128));
	wire w148128;
	torch #(1'b1) c148128 (.i_clk(tick), .i_in(), .o_out(w148128));
	wire w152128;
	torch #(1'b1) c152128 (.i_clk(tick), .i_in(), .o_out(w152128));
	wire w156128;
	torch #(1'b1) c156128 (.i_clk(tick), .i_in(), .o_out(w156128));
	wire w160128;
	torch #(1'b1) c160128 (.i_clk(tick), .i_in(), .o_out(w160128));
	wire w138131;
	repeater #(1, 1'b0, 0, 0) c138131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138131));
	wire w142131;
	repeater #(1, 1'b0, 0, 0) c142131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142131));
	wire w146131;
	repeater #(1, 1'b1, 0, 0) c146131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146131));
	wire w150131;
	repeater #(1, 1'b1, 0, 0) c150131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150131));
	wire w154131;
	repeater #(1, 1'b1, 0, 0) c154131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154131));
	wire w158131;
	repeater #(1, 1'b0, 0, 0) c158131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158131));
	wire w162131;
	repeater #(1, 1'b0, 0, 0) c162131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162131));
	wire w137132;
	repeater #(1, 1'b0, 0, 0) c137132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137132));
	wire w141132;
	repeater #(1, 1'b0, 0, 0) c141132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141132));
	wire w145132;
	repeater #(1, 1'b1, 0, 0) c145132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145132));
	wire w149132;
	repeater #(1, 1'b1, 0, 0) c149132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149132));
	wire w153132;
	repeater #(1, 1'b1, 0, 0) c153132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153132));
	wire w157132;
	repeater #(1, 1'b0, 0, 0) c157132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157132));
	wire w161132;
	repeater #(1, 1'b0, 0, 0) c161132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161132));
	wire w168132;
	repeater #(1, 1'b1, 0, 0) c168132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168132));
	wire w137166;
	torch #(1'b1) c137166 (.i_clk(tick), .i_in(), .o_out(w137166));
	wire w141166;
	torch #(1'b1) c141166 (.i_clk(tick), .i_in(), .o_out(w141166));
	wire w145166;
	torch #(1'b0) c145166 (.i_clk(tick), .i_in(), .o_out(w145166));
	wire w149166;
	torch #(1'b0) c149166 (.i_clk(tick), .i_in(), .o_out(w149166));
	wire w153166;
	torch #(1'b0) c153166 (.i_clk(tick), .i_in(), .o_out(w153166));
	wire w157166;
	torch #(1'b1) c157166 (.i_clk(tick), .i_in(), .o_out(w157166));
	wire w161166;
	torch #(1'b1) c161166 (.i_clk(tick), .i_in(), .o_out(w161166));
	wire w45171;

	wire w79171;

	wire w113171;

	wire w147171;

	wire w44172;
	repeater #(1, 1'b1, 0, 0) c44172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44172));
	wire w78172;
	repeater #(1, 1'b1, 0, 0) c78172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78172));
	wire w112172;
	repeater #(1, 1'b1, 0, 0) c112172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112172));
	wire w146172;
	repeater #(1, 1'b1, 0, 0) c146172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146172));
	wire w43173;

	wire w77173;

	wire w111173;

	wire w145173;

	wire w42174;
	repeater #(1, 1'b1, 0, 0) c42174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42174));
	wire w76174;
	repeater #(1, 1'b1, 0, 0) c76174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76174));
	wire w110174;
	repeater #(1, 1'b1, 0, 0) c110174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110174));
	wire w144174;
	repeater #(1, 1'b1, 0, 0) c144174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144174));
	wire w41175;

	wire w75175;

	wire w109175;

	wire w143175;

	wire w40176;
	repeater #(1, 1'b1, 0, 0) c40176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40176));
	wire w74176;
	repeater #(1, 1'b1, 0, 0) c74176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74176));
	wire w108176;
	repeater #(1, 1'b1, 0, 0) c108176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108176));
	wire w142176;
	repeater #(1, 1'b1, 0, 0) c142176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142176));
	wire w39177;

	wire w73177;

	wire w107177;

	wire w141177;

	wire w38178;
	repeater #(1, 1'b1, 0, 0) c38178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38178));
	wire w72178;
	repeater #(1, 1'b1, 0, 0) c72178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72178));
	wire w106178;
	repeater #(1, 1'b1, 0, 0) c106178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106178));
	wire w140178;
	repeater #(1, 1'b1, 0, 0) c140178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140178));
	wire w37179;

	wire w71179;

	wire w105179;

	wire w139179;

	wire w36180;
	repeater #(1, 1'b0, 0, 0) c36180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36180));
	wire w70180;
	repeater #(1, 1'b0, 0, 0) c70180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70180));
	wire w104180;
	repeater #(1, 1'b0, 0, 0) c104180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104180));
	wire w138180;
	repeater #(1, 1'b0, 0, 0) c138180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138180));
	wire w35181;

	wire w69181;

	wire w103181;

	wire w137181;

	wire w34182;
	repeater #(1, 1'b0, 0, 0) c34182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34182));
	wire w68182;
	repeater #(1, 1'b0, 0, 0) c68182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68182));
	wire w102182;
	repeater #(1, 1'b0, 0, 0) c102182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102182));
	wire w136182;
	repeater #(1, 1'b0, 0, 0) c136182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136182));
	wire w33183;

	wire w67183;

	wire w101183;

	wire w135183;

	wire w32184;
	repeater #(1, 1'b1, 0, 0) c32184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32184));
	wire w66184;
	repeater #(1, 1'b1, 0, 0) c66184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66184));
	wire w100184;
	repeater #(1, 1'b1, 0, 0) c100184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100184));
	wire w134184;
	repeater #(1, 1'b1, 0, 0) c134184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134184));
	wire w31185;

	wire w65185;

	wire w99185;

	wire w133185;

	wire w30186;
	repeater #(1, 1'b0, 0, 0) c30186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30186));
	wire w64186;
	repeater #(1, 1'b0, 0, 0) c64186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64186));
	wire w98186;
	repeater #(1, 1'b0, 0, 0) c98186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98186));
	wire w132186;
	repeater #(1, 1'b0, 0, 0) c132186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132186));
	wire w29187;

	wire w63187;

	wire w97187;

	wire w131187;

	wire w28188;
	repeater #(1, 1'b0, 0, 0) c28188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28188));
	wire w62188;
	repeater #(1, 1'b0, 0, 0) c62188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62188));
	wire w96188;
	repeater #(1, 1'b0, 0, 0) c96188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96188));
	wire w130188;
	repeater #(1, 1'b0, 0, 0) c130188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130188));
	wire w27189;

	wire w61189;

	wire w95189;

	wire w129189;

	wire w26190;
	repeater #(1, 1'b0, 0, 0) c26190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26190));
	wire w60190;
	repeater #(1, 1'b0, 0, 0) c60190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60190));
	wire w94190;
	repeater #(1, 1'b0, 0, 0) c94190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94190));
	wire w128190;
	repeater #(1, 1'b0, 0, 0) c128190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128190));
	wire w25191;

	wire w59191;

	wire w93191;

	wire w127191;

	wire w24192;
	repeater #(1, 1'b1, 0, 0) c24192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24192));
	wire w58192;
	repeater #(1, 1'b1, 0, 0) c58192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58192));
	wire w92192;
	repeater #(1, 1'b1, 0, 0) c92192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92192));
	wire w126192;
	repeater #(1, 1'b1, 0, 0) c126192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126192));
	wire w23193;

	wire w57193;

	wire w91193;

	wire w125193;

	wire w22194;
	repeater #(1, 1'b1, 0, 0) c22194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22194));
	wire w56194;
	repeater #(1, 1'b1, 0, 0) c56194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56194));
	wire w90194;
	repeater #(1, 1'b1, 0, 0) c90194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90194));
	wire w124194;
	repeater #(1, 1'b1, 0, 0) c124194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124194));
	wire w21195;

	wire w55195;

	wire w89195;

	wire w123195;

	wire w20196;
	repeater #(1, 1'b1, 0, 0) c20196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20196));
	wire w54196;
	repeater #(1, 1'b1, 0, 0) c54196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54196));
	wire w88196;
	repeater #(1, 1'b1, 0, 0) c88196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88196));
	wire w122196;
	repeater #(1, 1'b1, 0, 0) c122196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122196));
	wire w19197;

	wire w53197;

	wire w87197;

	wire w121197;

	wire w18198;
	repeater #(1, 1'b1, 0, 0) c18198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18198));
	wire w52198;
	repeater #(1, 1'b1, 0, 0) c52198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52198));
	wire w86198;
	repeater #(1, 1'b1, 0, 0) c86198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86198));
	wire w120198;
	repeater #(1, 1'b1, 0, 0) c120198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120198));
	wire w161103;
	repeater #(2, 1'b1, 0, 0) c161103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161103));
	wire w501103;
	repeater #(2, 1'b1, 0, 0) c501103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w501103));
	wire w1361104;
	repeater #(1, 1'b1, 0, 0) c1361104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361104));
	wire w1401104;
	repeater #(1, 1'b1, 0, 0) c1401104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401104));
	wire w1441104;
	repeater #(1, 1'b0, 0, 0) c1441104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441104));
	wire w1481104;
	repeater #(1, 1'b0, 0, 0) c1481104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1481104));
	wire w1521104;
	repeater #(1, 1'b0, 0, 0) c1521104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1521104));
	wire w1561104;
	repeater #(1, 1'b1, 0, 0) c1561104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1561104));
	wire w1601104;
	repeater #(1, 1'b1, 0, 0) c1601104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1601104));
	wire w21105;
	repeater #(1, 1'b1, 0, 0) c21105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21105));
	wire w81105;
	torch #(1'b1) c81105 (.i_clk(tick), .i_in(), .o_out(w81105));
	wire w181105;
	repeater #(1, 1'b1, 0, 0) c181105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181105));
	wire w241105;
	torch #(1'b1) c241105 (.i_clk(tick), .i_in(), .o_out(w241105));
	wire w361105;
	repeater #(1, 1'b1, 0, 0) c361105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w361105));
	wire w421105;
	torch #(1'b1) c421105 (.i_clk(tick), .i_in(), .o_out(w421105));
	wire w521105;
	repeater #(1, 1'b1, 0, 0) c521105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w521105));
	wire w581105;
	torch #(1'b1) c581105 (.i_clk(tick), .i_in(), .o_out(w581105));
	wire w1361105;
	repeater #(1, 1'b1, 0, 0) c1361105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361105));
	wire w1381105;
	repeater #(1, 1'b0, 0, 0) c1381105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1381105));
	wire w1401105;
	repeater #(1, 1'b1, 0, 0) c1401105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401105));
	wire w1421105;
	repeater #(1, 1'b0, 0, 0) c1421105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1421105));
	wire w1441105;
	repeater #(1, 1'b0, 0, 0) c1441105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441105));
	wire w1461105;
	repeater #(1, 1'b0, 0, 0) c1461105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1461105));
	wire w1481105;
	repeater #(1, 1'b0, 0, 0) c1481105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1481105));
	wire w1501105;
	repeater #(1, 1'b0, 0, 0) c1501105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1501105));
	wire w1521105;
	repeater #(1, 1'b0, 0, 0) c1521105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1521105));
	wire w1541105;
	repeater #(1, 1'b0, 0, 0) c1541105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541105));
	wire w1561105;
	repeater #(1, 1'b1, 0, 0) c1561105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1561105));
	wire w1581105;
	repeater #(1, 1'b0, 0, 0) c1581105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581105));
	wire w1601105;
	repeater #(1, 1'b1, 0, 0) c1601105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1601105));
	wire w1621105;
	repeater #(1, 1'b0, 0, 0) c1621105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621105));
	wire w1371106;
	torch #(1'b0) c1371106 (.i_clk(tick), .i_in(), .o_out(w1371106));
	wire w1411106;
	torch #(1'b0) c1411106 (.i_clk(tick), .i_in(), .o_out(w1411106));
	wire w1451106;
	torch #(1'b0) c1451106 (.i_clk(tick), .i_in(), .o_out(w1451106));
	wire w1491106;
	torch #(1'b0) c1491106 (.i_clk(tick), .i_in(), .o_out(w1491106));
	wire w1531106;
	torch #(1'b0) c1531106 (.i_clk(tick), .i_in(), .o_out(w1531106));
	wire w1571106;
	torch #(1'b0) c1571106 (.i_clk(tick), .i_in(), .o_out(w1571106));
	wire w1611106;
	torch #(1'b0) c1611106 (.i_clk(tick), .i_in(), .o_out(w1611106));
	wire w91108;
	repeater #(1, 1'b1, 0, 0) c91108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91108));
	wire w431108;
	repeater #(1, 1'b1, 0, 0) c431108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w431108));
	wire w21109;
	repeater #(1, 1'b1, 0, 0) c21109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21109));
	wire w181109;
	repeater #(1, 1'b1, 0, 0) c181109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181109));
	wire w361109;
	repeater #(1, 1'b1, 0, 0) c361109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w361109));
	wire w521109;
	repeater #(1, 1'b1, 0, 0) c521109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w521109));
	wire w771109;
	repeater #(1, 1'b1, 0, 0) c771109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w771109));
	wire w811109;
	repeater #(1, 1'b1, 0, 0) c811109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811109));
	wire w851109;
	repeater #(1, 1'b1, 0, 0) c851109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w851109));
	wire w891109;
	repeater #(1, 1'b1, 0, 0) c891109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w891109));
	wire w1091109;
	repeater #(1, 1'b0, 0, 0) c1091109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1091109));
	wire w1131109;
	repeater #(1, 1'b0, 0, 0) c1131109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1131109));
	wire w1171109;
	repeater #(1, 1'b0, 0, 0) c1171109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171109));
	wire w1211109;
	repeater #(1, 1'b0, 0, 0) c1211109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1211109));
	wire w71110;

	wire w231110;

	wire w411110;

	wire w571110;

	wire w151111;

	wire w491111;

	wire w11112;

	wire w21112;

	wire w121112;

	wire w171112;

	wire w181112;

	wire w351112;

	wire w361112;

	wire w461112;

	wire w511112;

	wire w521112;

	wire w101114;

	wire w441114;

	wire w01115;

	wire w11115;

	wire w161115;

	wire w171115;

	wire w341115;

	wire w351115;

	wire w501115;

	wire w511115;

	wire w21116;

	wire w61116;

	wire w101116;

	wire w361116;

	wire w401116;

	wire w441116;

	wire w1381116;

	wire w1421116;

	wire w1461116;

	wire w1501116;

	wire w1541116;

	wire w1581116;

	wire w1621116;

	wire w261119;

	wire w601119;

	wire w2071119;

	wire w01120;

	wire w31120;

	wire w41120;

	wire w71120;

	wire w81120;

	wire w111120;

	wire w121120;

	wire w151120;

	wire w161120;

	wire w191120;

	wire w201120;

	wire w231120;

	wire w241120;

	wire w331120;

	wire w341120;

	wire w371120;

	wire w381120;

	wire w411120;

	wire w421120;

	wire w451120;

	wire w461120;

	wire w491120;

	wire w501120;

	wire w531120;

	wire w541120;

	wire w571120;

	wire w581120;

	wire w2051120;

	wire w311121;

	wire w821123;

	wire w851123;

	wire w1131123;

	wire w1161123;

	wire w121124;
	repeater #(1, 1'b1, 0, 0) c121124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121124));
	wire w161124;
	repeater #(1, 1'b1, 0, 0) c161124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161124));
	wire w201124;
	repeater #(1, 1'b1, 0, 0) c201124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201124));
	wire w461124;
	repeater #(1, 1'b1, 0, 0) c461124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w461124));
	wire w501124;
	repeater #(1, 1'b1, 0, 0) c501124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w501124));
	wire w541124;
	repeater #(1, 1'b1, 0, 0) c541124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w541124));
	wire w711126;
	repeater #(1, 1'b1, 0, 0) c711126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711126));
	wire w761126;
	repeater #(1, 1'b1, 0, 0) c761126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761126));
	wire w811126;
	repeater #(1, 1'b1, 0, 0) c811126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811126));
	wire w1171126;
	repeater #(1, 1'b0, 0, 0) c1171126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171126));
	wire w1221126;
	repeater #(1, 1'b1, 0, 0) c1221126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221126));
	wire w1271126;
	repeater #(1, 1'b1, 0, 0) c1271126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271126));
	wire w2061126;

	wire w21127;

	wire w181127;

	wire w221127;

	wire w321127;

	wire w361127;

	wire w521127;

	wire w561127;

	wire w701127;

	wire w711127;
	repeater #(1, 1'b1, 0, 0) c711127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711127));
	wire w751127;

	wire w761127;
	repeater #(1, 1'b1, 0, 0) c761127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761127));
	wire w801127;

	wire w811127;
	repeater #(1, 1'b1, 0, 0) c811127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811127));
	wire w1171127;
	repeater #(1, 1'b0, 0, 0) c1171127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171127));
	wire w1181127;

	wire w1221127;
	repeater #(1, 1'b1, 0, 0) c1221127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221127));
	wire w1231127;

	wire w1271127;
	repeater #(1, 1'b1, 0, 0) c1271127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271127));
	wire w1281127;

	wire w1381127;
	torch #(1'b0) c1381127 (.i_clk(tick), .i_in(), .o_out(w1381127));
	wire w1421127;
	torch #(1'b0) c1421127 (.i_clk(tick), .i_in(), .o_out(w1421127));
	wire w1461127;
	torch #(1'b1) c1461127 (.i_clk(tick), .i_in(), .o_out(w1461127));
	wire w1501127;
	torch #(1'b1) c1501127 (.i_clk(tick), .i_in(), .o_out(w1501127));
	wire w1541127;
	torch #(1'b1) c1541127 (.i_clk(tick), .i_in(), .o_out(w1541127));
	wire w1581127;
	torch #(1'b0) c1581127 (.i_clk(tick), .i_in(), .o_out(w1581127));
	wire w1621127;
	torch #(1'b0) c1621127 (.i_clk(tick), .i_in(), .o_out(w1621127));
	wire w01128;
	repeater #(1, 1'b1, 0, 0) c01128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w01128));
	wire w161128;
	repeater #(1, 1'b1, 0, 0) c161128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161128));
	wire w341128;
	repeater #(1, 1'b1, 0, 0) c341128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w341128));
	wire w501128;
	repeater #(1, 1'b1, 0, 0) c501128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w501128));
	wire w71129;
	repeater #(1, 1'b1, 0, 0) c71129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71129));
	wire w411129;
	repeater #(1, 1'b0, 0, 0) c411129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w411129));
	wire w21130;

	wire w181130;

	wire w361130;

	wire w521130;

	wire w711130;
	repeater #(1, 1'b1, 0, 0) c711130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711130));
	wire w761130;
	repeater #(1, 1'b0, 0, 0) c761130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761130));
	wire w811130;
	repeater #(1, 1'b0, 0, 0) c811130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811130));
	wire w1171130;
	repeater #(1, 1'b0, 0, 0) c1171130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171130));
	wire w1221130;
	repeater #(1, 1'b1, 0, 0) c1221130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221130));
	wire w1271130;
	repeater #(1, 1'b1, 0, 0) c1271130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271130));
	wire w101131;

	wire w441131;

	wire w701131;

	wire w711131;
	repeater #(1, 1'b0, 0, 0) c711131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711131));
	wire w751131;

	wire w761131;
	repeater #(1, 1'b0, 0, 0) c761131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761131));
	wire w801131;

	wire w811131;
	repeater #(1, 1'b0, 0, 0) c811131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811131));
	wire w1171131;
	repeater #(1, 1'b0, 0, 0) c1171131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171131));
	wire w1181131;

	wire w1221131;
	repeater #(1, 1'b1, 0, 0) c1221131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221131));
	wire w1231131;

	wire w1271131;
	repeater #(1, 1'b1, 0, 0) c1271131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271131));
	wire w1281131;

	wire w51132;

	wire w71132;

	wire w81132;

	wire w131132;

	wire w211132;

	wire w391132;

	wire w411132;

	wire w421132;

	wire w471132;

	wire w551132;

	wire w1381132;

	wire w1421132;

	wire w1461132;

	wire w1501132;

	wire w1541132;

	wire w1581132;

	wire w1621132;

	wire w151134;

	wire w161134;

	wire w491134;

	wire w501134;

	wire w711134;
	repeater #(1, 1'b0, 0, 0) c711134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711134));
	wire w761134;
	repeater #(1, 1'b0, 0, 0) c761134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761134));
	wire w811134;
	repeater #(1, 1'b0, 0, 0) c811134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811134));
	wire w1171134;
	repeater #(1, 1'b0, 0, 0) c1171134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171134));
	wire w1221134;
	repeater #(1, 1'b1, 0, 0) c1221134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221134));
	wire w1271134;
	repeater #(1, 1'b1, 0, 0) c1271134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271134));
	wire w701135;

	wire w711135;
	repeater #(1, 1'b0, 0, 0) c711135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711135));
	wire w751135;

	wire w761135;
	repeater #(1, 1'b0, 0, 0) c761135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761135));
	wire w801135;

	wire w811135;
	repeater #(1, 1'b0, 0, 0) c811135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w811135));
	wire w1171135;
	repeater #(1, 1'b0, 0, 0) c1171135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171135));
	wire w1181135;

	wire w1221135;
	repeater #(1, 1'b1, 0, 0) c1221135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221135));
	wire w1231135;

	wire w1271135;
	repeater #(1, 1'b1, 0, 0) c1271135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271135));
	wire w1281135;

	wire w51136;

	wire w71136;

	wire w81136;

	wire w500;

	wire w2300;

	wire w2500;

	wire w2600;

	wire w3900;

	wire w19401;
	torch #(1'b1) c19401 (.i_clk(tick), .i_in(), .o_out(w19401));
	wire w19501;

	wire w202;
	torch #(1'b1) c202 (.i_clk(tick), .i_in(), .o_out(w202));
	wire w302;

	wire w2002;
	torch #(1'b1) c2002 (.i_clk(tick), .i_in(), .o_out(w2002));
	wire w2102;

	wire w3602;
	torch #(1'b1) c3602 (.i_clk(tick), .i_in(), .o_out(w3602));
	wire w3702;

	wire w5602;
	repeater #(2, 1'b1, 0, 0) c5602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5602));
	wire w11002;
	repeater #(2, 1'b1, 0, 0) c11002 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11002));
	wire w19502;

	wire w19702;

	wire w303;

	wire w503;

	wire w2103;

	wire w2303;

	wire w3703;

	wire w3903;

	wire w5303;
	repeater #(1, 1'b1, 0, 0) c5303 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5303));
	wire w6103;
	repeater #(1, 1'b0, 0, 0) c6103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6103));
	wire w6203;
	repeater #(2, 1'b0, 0, 0) c6203 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6203));
	wire w10403;
	repeater #(2, 1'b0, 0, 0) c10403 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10403));
	wire w10503;
	repeater #(1, 1'b0, 0, 0) c10503 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10503));
	wire w11303;
	repeater #(1, 1'b1, 0, 0) c11303 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11303));
	wire w5704;
	repeater #(1, 1'b0, 0, 0) c5704 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5704));
	wire w10904;
	repeater #(1, 1'b0, 0, 0) c10904 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10904));
	wire w19704;

	wire w19804;

	wire w19904;

	wire w505;

	wire w605;

	wire w705;

	wire w2305;

	wire w2405;

	wire w2505;

	wire w3905;

	wire w4005;

	wire w4105;

	wire w6305;

	wire w6705;
	repeater #(1, 1'b0, 0, 0) c6705 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6705));
	wire w9905;
	repeater #(1, 1'b1, 0, 0) c9905 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9905));
	wire w10305;

	wire w19205;

	wire w19305;

	wire w19905;

	wire w006;

	wire w106;

	wire w706;

	wire w1806;

	wire w1906;

	wire w2506;

	wire w3406;

	wire w3506;

	wire w4106;

	wire w6406;

	wire w10206;

	wire w6307;
	repeater #(2, 1'b0, 0, 0) c6307 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6307));
	wire w10307;
	repeater #(2, 1'b1, 0, 0) c10307 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10307));
	wire w12207;
	torch #(1'b0) c12207 (.i_clk(tick), .i_in(), .o_out(w12207));
	wire w12607;
	torch #(1'b0) c12607 (.i_clk(tick), .i_in(), .o_out(w12607));
	wire w13007;
	torch #(1'b1) c13007 (.i_clk(tick), .i_in(), .o_out(w13007));
	wire w13407;
	torch #(1'b1) c13407 (.i_clk(tick), .i_in(), .o_out(w13407));
	wire w13807;
	torch #(1'b1) c13807 (.i_clk(tick), .i_in(), .o_out(w13807));
	wire w14207;
	torch #(1'b0) c14207 (.i_clk(tick), .i_in(), .o_out(w14207));
	wire w14607;
	torch #(1'b0) c14607 (.i_clk(tick), .i_in(), .o_out(w14607));
	wire w19707;
	repeater #(1, 1'b0, 0, 0) c19707 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19707));
	wire w19907;
	torch #(1'b0) c19907 (.i_clk(tick), .i_in(), .o_out(w19907));
	wire w20507;
	torch #(1'b1) c20507 (.i_clk(tick), .i_in(), .o_out(w20507));
	wire w508;
	repeater #(1, 1'b0, 0, 0) c508 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w508));
	wire w708;
	torch #(1'b0) c708 (.i_clk(tick), .i_in(), .o_out(w708));
	wire w2308;
	repeater #(1, 1'b0, 0, 0) c2308 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2308));
	wire w2508;
	torch #(1'b0) c2508 (.i_clk(tick), .i_in(), .o_out(w2508));
	wire w3108;
	torch #(1'b1) c3108 (.i_clk(tick), .i_in(), .o_out(w3108));
	wire w3908;
	repeater #(1, 1'b0, 0, 0) c3908 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3908));
	wire w4108;
	torch #(1'b0) c4108 (.i_clk(tick), .i_in(), .o_out(w4108));
	wire w5708;

	wire w5808;

	wire w10808;

	wire w10908;

	wire w5609;

	wire w6509;

	wire w10109;

	wire w11009;

	wire w20109;
	repeater #(1, 1'b1, 0, 0) c20109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20109));
	wire w9010;
	repeater #(1, 1'b1, 0, 0) c9010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9010));
	wire w27010;
	repeater #(1, 1'b1, 0, 0) c27010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27010));
	wire w43010;
	repeater #(1, 1'b1, 0, 0) c43010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43010));
	wire w59010;

	wire w107010;

	wire w198011;
	torch #(1'b1) c198011 (.i_clk(tick), .i_in(), .o_out(w198011));
	wire w6012;
	torch #(1'b1) c6012 (.i_clk(tick), .i_in(), .o_out(w6012));
	wire w24012;
	torch #(1'b1) c24012 (.i_clk(tick), .i_in(), .o_out(w24012));
	wire w40012;
	torch #(1'b1) c40012 (.i_clk(tick), .i_in(), .o_out(w40012));
	wire w122012;

	wire w126012;

	wire w130012;

	wire w134012;

	wire w138012;

	wire w142012;

	wire w146012;

	wire w206013;
	torch #(1'b1) c206013 (.i_clk(tick), .i_in(), .o_out(w206013));
	wire w32014;
	torch #(1'b1) c32014 (.i_clk(tick), .i_in(), .o_out(w32014));
	wire w197014;
	repeater #(1, 1'b0, 0, 0) c197014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197014));
	wire w5015;
	repeater #(1, 1'b0, 0, 0) c5015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5015));
	wire w23015;
	repeater #(1, 1'b0, 0, 0) c23015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23015));
	wire w39015;
	repeater #(1, 1'b0, 0, 0) c39015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39015));
	wire w207015;
	repeater #(1, 1'b0, 0, 0) c207015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207015));
	wire w11016;
	repeater #(1, 1'b0, 0, 0) c11016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11016));
	wire w33016;
	repeater #(1, 1'b0, 0, 0) c33016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33016));
	wire w45016;
	repeater #(1, 1'b0, 0, 0) c45016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45016));
	wire w11018;
	repeater #(1, 1'b0, 0, 0) c11018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11018));
	wire w45018;
	repeater #(1, 1'b0, 0, 0) c45018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45018));
	wire w122023;
	torch #(1'b0) c122023 (.i_clk(tick), .i_in(), .o_out(w122023));
	wire w126023;
	torch #(1'b0) c126023 (.i_clk(tick), .i_in(), .o_out(w126023));
	wire w130023;
	torch #(1'b1) c130023 (.i_clk(tick), .i_in(), .o_out(w130023));
	wire w134023;
	torch #(1'b1) c134023 (.i_clk(tick), .i_in(), .o_out(w134023));
	wire w138023;
	torch #(1'b1) c138023 (.i_clk(tick), .i_in(), .o_out(w138023));
	wire w142023;
	torch #(1'b0) c142023 (.i_clk(tick), .i_in(), .o_out(w142023));
	wire w146023;
	torch #(1'b0) c146023 (.i_clk(tick), .i_in(), .o_out(w146023));
	wire w122028;

	wire w126028;

	wire w130028;

	wire w134028;

	wire w138028;

	wire w142028;

	wire w146028;

	wire w122039;
	torch #(1'b0) c122039 (.i_clk(tick), .i_in(), .o_out(w122039));
	wire w126039;
	torch #(1'b0) c126039 (.i_clk(tick), .i_in(), .o_out(w126039));
	wire w130039;
	torch #(1'b1) c130039 (.i_clk(tick), .i_in(), .o_out(w130039));
	wire w134039;
	torch #(1'b1) c134039 (.i_clk(tick), .i_in(), .o_out(w134039));
	wire w138039;
	torch #(1'b1) c138039 (.i_clk(tick), .i_in(), .o_out(w138039));
	wire w142039;
	torch #(1'b0) c142039 (.i_clk(tick), .i_in(), .o_out(w142039));
	wire w146039;
	torch #(1'b0) c146039 (.i_clk(tick), .i_in(), .o_out(w146039));
	wire w122044;

	wire w126044;

	wire w130044;

	wire w134044;

	wire w138044;

	wire w142044;

	wire w146044;

	wire w122055;
	torch #(1'b0) c122055 (.i_clk(tick), .i_in(), .o_out(w122055));
	wire w126055;
	torch #(1'b0) c126055 (.i_clk(tick), .i_in(), .o_out(w126055));
	wire w130055;
	torch #(1'b1) c130055 (.i_clk(tick), .i_in(), .o_out(w130055));
	wire w134055;
	torch #(1'b1) c134055 (.i_clk(tick), .i_in(), .o_out(w134055));
	wire w138055;
	torch #(1'b1) c138055 (.i_clk(tick), .i_in(), .o_out(w138055));
	wire w142055;
	torch #(1'b0) c142055 (.i_clk(tick), .i_in(), .o_out(w142055));
	wire w146055;
	torch #(1'b0) c146055 (.i_clk(tick), .i_in(), .o_out(w146055));
	wire w120058;
	assign outputs[1] = ();
	wire w122058;
	assign outputs[2] = ();
	wire w124058;
	assign outputs[3] = ();
	wire w126058;
	assign outputs[4] = ();
	wire w128058;
	assign outputs[5] = ();
	wire w130058;
	assign outputs[6] = ();
	wire w132058;
	assign outputs[7] = ();
	wire w134058;
	assign outputs[8] = ();
	wire w136058;
	assign outputs[9] = ();
	wire w138058;
	assign outputs[10] = ();
	wire w140058;
	assign outputs[11] = ();
	wire w142058;
	assign outputs[12] = ();
	wire w144058;
	assign outputs[13] = ();
	wire w146058;
	assign outputs[14] = ();
	wire w120059;
	repeater #(1, 1'b0, 0, 0) c120059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120059));
	wire w122059;
	repeater #(1, 1'b0, 0, 0) c122059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122059));
	wire w124059;
	repeater #(1, 1'b0, 0, 0) c124059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124059));
	wire w126059;
	repeater #(1, 1'b0, 0, 0) c126059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126059));
	wire w128059;
	repeater #(1, 1'b1, 0, 0) c128059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128059));
	wire w130059;
	repeater #(1, 1'b1, 0, 0) c130059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130059));
	wire w132059;
	repeater #(1, 1'b0, 0, 0) c132059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132059));
	wire w134059;
	repeater #(1, 1'b1, 0, 0) c134059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134059));
	wire w136059;
	repeater #(1, 1'b1, 0, 0) c136059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136059));
	wire w138059;
	repeater #(1, 1'b1, 0, 0) c138059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138059));
	wire w140059;
	repeater #(1, 1'b0, 0, 0) c140059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140059));
	wire w142059;
	repeater #(1, 1'b0, 0, 0) c142059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142059));
	wire w144059;
	repeater #(1, 1'b0, 0, 0) c144059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144059));
	wire w146059;
	repeater #(1, 1'b0, 0, 0) c146059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146059));
	wire w121066;
	repeater #(2, 1'b1, 0, 0) c121066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121066));
	wire w125066;
	repeater #(2, 1'b1, 0, 0) c125066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125066));
	wire w129066;
	repeater #(2, 1'b0, 0, 0) c129066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w129066));
	wire w133066;
	repeater #(2, 1'b0, 0, 0) c133066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133066));
	wire w137066;
	repeater #(2, 1'b0, 0, 0) c137066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137066));
	wire w141066;
	repeater #(2, 1'b1, 0, 0) c141066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141066));
	wire w145066;
	repeater #(2, 1'b1, 0, 0) c145066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145066));
	wire w119071;
	repeater #(1, 1'b1, 0, 0) c119071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119071));
	wire w121071;
	assign w121071 = inputs[6];
	wire w123071;
	repeater #(1, 1'b1, 0, 0) c123071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123071));
	wire w125071;
	assign w125071 = inputs[7];
	wire w127071;
	repeater #(1, 1'b0, 0, 0) c127071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127071));
	wire w129071;
	assign w129071 = inputs[8];
	wire w131071;
	repeater #(1, 1'b0, 0, 0) c131071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131071));
	wire w133071;
	assign w133071 = inputs[9];
	wire w135071;
	repeater #(1, 1'b0, 0, 0) c135071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135071));
	wire w137071;
	assign w137071 = inputs[10];
	wire w139071;
	repeater #(1, 1'b1, 0, 0) c139071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139071));
	wire w143071;
	repeater #(1, 1'b1, 0, 0) c143071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143071));
	wire w145071;
	assign w145071 = inputs[11];
	wire w121072;

	wire w125072;

	wire w129072;

	wire w133072;

	wire w137072;

	wire w141072;

	wire w145072;

	wire w120073;

	wire w124073;

	wire w128073;

	wire w132073;

	wire w136073;

	wire w140073;

	wire w144073;

	wire w121074;
	torch #(1'b1) c121074 (.i_clk(tick), .i_in(), .o_out(w121074));
	wire w125074;
	torch #(1'b1) c125074 (.i_clk(tick), .i_in(), .o_out(w125074));
	wire w129074;
	torch #(1'b1) c129074 (.i_clk(tick), .i_in(), .o_out(w129074));
	wire w133074;
	torch #(1'b1) c133074 (.i_clk(tick), .i_in(), .o_out(w133074));
	wire w137074;
	torch #(1'b1) c137074 (.i_clk(tick), .i_in(), .o_out(w137074));
	wire w141074;
	torch #(1'b1) c141074 (.i_clk(tick), .i_in(), .o_out(w141074));
	wire w145074;
	torch #(1'b1) c145074 (.i_clk(tick), .i_in(), .o_out(w145074));
	wire w119075;
	repeater #(1, 1'b1, 0, 0) c119075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119075));
	wire w123075;
	repeater #(1, 1'b1, 0, 0) c123075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123075));
	wire w127075;
	repeater #(1, 1'b1, 0, 0) c127075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127075));
	wire w131075;
	repeater #(1, 1'b1, 0, 0) c131075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131075));
	wire w135075;
	repeater #(1, 1'b1, 0, 0) c135075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135075));
	wire w139075;
	repeater #(1, 1'b1, 0, 0) c139075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139075));
	wire w143075;
	repeater #(1, 1'b1, 0, 0) c143075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143075));
	wire w1460133;

	wire w1440135;

	wire w1420137;

	wire w1400139;

	wire w1380141;

	wire w2040145;
	repeater #(2, 1'b0, 0, 0) c2040145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040145));
	wire w300146;
	repeater #(2, 1'b0, 0, 0) c300146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300146));
	wire w1210147;
	torch #(1'b1) c1210147 (.i_clk(tick), .i_in(), .o_out(w1210147));
	wire w1250147;
	torch #(1'b1) c1250147 (.i_clk(tick), .i_in(), .o_out(w1250147));
	wire w1290147;
	torch #(1'b1) c1290147 (.i_clk(tick), .i_in(), .o_out(w1290147));
	wire w1330147;
	torch #(1'b1) c1330147 (.i_clk(tick), .i_in(), .o_out(w1330147));
	wire w1370147;
	torch #(1'b1) c1370147 (.i_clk(tick), .i_in(), .o_out(w1370147));
	wire w1410147;
	torch #(1'b1) c1410147 (.i_clk(tick), .i_in(), .o_out(w1410147));
	wire w1450147;
	torch #(1'b1) c1450147 (.i_clk(tick), .i_in(), .o_out(w1450147));
	wire w1960147;
	torch #(1'b1) c1960147 (.i_clk(tick), .i_in(), .o_out(w1960147));
	wire w2060147;
	repeater #(1, 1'b1, 0, 0) c2060147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060147));
	wire w40148;
	torch #(1'b1) c40148 (.i_clk(tick), .i_in(), .o_out(w40148));
	wire w220148;
	torch #(1'b1) c220148 (.i_clk(tick), .i_in(), .o_out(w220148));
	wire w320148;
	repeater #(1, 1'b0, 0, 0) c320148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320148));
	wire w380148;
	torch #(1'b1) c380148 (.i_clk(tick), .i_in(), .o_out(w380148));
	wire w1220150;
	repeater #(2, 1'b0, 0, 0) c1220150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1220150));
	wire w1260150;
	repeater #(2, 1'b0, 0, 0) c1260150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1260150));
	wire w1300150;
	repeater #(2, 1'b0, 0, 0) c1300150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1300150));
	wire w1340150;
	repeater #(2, 1'b0, 0, 0) c1340150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340150));
	wire w1380150;
	repeater #(1, 1'b0, 0, 0) c1380150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380150));
	wire w1420150;
	repeater #(1, 1'b0, 0, 0) c1420150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420150));
	wire w1460150;
	repeater #(1, 1'b0, 0, 0) c1460150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460150));
	wire w1970150;
	repeater #(1, 1'b1, 0, 0) c1970150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970150));
	wire w50151;
	repeater #(1, 1'b1, 0, 0) c50151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50151));
	wire w230151;
	repeater #(1, 1'b1, 0, 0) c230151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230151));
	wire w390151;
	repeater #(1, 1'b1, 0, 0) c390151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390151));
	wire w1350151;
	repeater #(1, 1'b0, 0, 0) c1350151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350151));
	wire w1470151;
	repeater #(2, 1'b0, 0, 0) c1470151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470151));
	wire w1490151;
	torch #(1'b1) c1490151 (.i_clk(tick), .i_in(), .o_out(w1490151));
	wire w2060151;
	repeater #(1, 1'b1, 0, 0) c2060151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060151));
	wire w320152;
	repeater #(1, 1'b0, 0, 0) c320152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320152));
	wire w1950152;

	wire w30153;

	wire w210153;

	wire w370153;

	wire w2030153;

	wire w290154;

	wire w2000154;

	wire w2050154;

	wire w2060154;

	wire w260155;

	wire w310155;

	wire w320155;

	wire w1240156;
	repeater #(1, 1'b0, 0, 0) c1240156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240156));
	wire w1440156;
	repeater #(1, 1'b0, 0, 0) c1440156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1440156));
	wire w1980156;

	wire w60157;

	wire w240157;

	wire w400157;

	wire w2040157;

	wire w2050157;

	wire w300158;

	wire w310158;

	wire w1900158;

	wire w160159;

	wire w590159;
	repeater #(2, 1'b0, 0, 0) c590159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590159));
	wire w610159;
	repeater #(1, 1'b1, 0, 0) c610159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w610159));
	wire w630159;
	repeater #(2, 1'b0, 0, 0) c630159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630159));
	wire w650159;
	repeater #(1, 1'b1, 0, 0) c650159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650159));
	wire w670159;
	repeater #(2, 1'b0, 0, 0) c670159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w670159));
	wire w690159;
	repeater #(1, 1'b1, 0, 0) c690159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w690159));
	wire w710159;
	repeater #(2, 1'b0, 0, 0) c710159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710159));
	wire w730159;
	repeater #(1, 1'b1, 0, 0) c730159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w730159));
	wire w930159;
	repeater #(1, 1'b0, 0, 0) c930159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w930159));
	wire w950159;
	repeater #(2, 1'b0, 0, 0) c950159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w950159));
	wire w970159;
	repeater #(1, 1'b0, 0, 0) c970159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w970159));
	wire w990159;
	repeater #(2, 1'b0, 0, 0) c990159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990159));
	wire w1010159;
	repeater #(1, 1'b0, 0, 0) c1010159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010159));
	wire w1030159;
	repeater #(2, 1'b0, 0, 0) c1030159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030159));
	wire w1050159;
	repeater #(1, 1'b0, 0, 0) c1050159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1050159));
	wire w1070159;
	repeater #(2, 1'b0, 0, 0) c1070159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070159));
	wire w1910160;
	repeater #(1, 1'b1, 0, 0) c1910160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910160));
	wire w1950160;
	repeater #(1, 1'b1, 0, 0) c1950160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950160));
	wire w1990160;
	repeater #(1, 1'b1, 0, 0) c1990160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990160));
	wire w2030160;
	repeater #(1, 1'b1, 0, 0) c2030160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030160));
	wire w2070160;
	repeater #(1, 1'b1, 0, 0) c2070160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070160));
	wire w30161;
	repeater #(1, 1'b1, 0, 0) c30161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30161));
	wire w70161;
	repeater #(1, 1'b1, 0, 0) c70161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70161));
	wire w170161;
	repeater #(1, 1'b1, 0, 0) c170161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170161));
	wire w210161;
	repeater #(1, 1'b1, 0, 0) c210161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210161));
	wire w250161;
	repeater #(1, 1'b1, 0, 0) c250161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250161));
	wire w290161;
	repeater #(1, 1'b0, 0, 0) c290161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290161));
	wire w330161;
	repeater #(1, 1'b1, 0, 0) c330161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330161));
	wire w370161;
	repeater #(1, 1'b1, 0, 0) c370161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370161));
	wire w410161;
	repeater #(1, 1'b1, 0, 0) c410161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w410161));
	wire w680161;

	wire w980161;

	wire w600162;

	wire w640162;

	wire w670162;

	wire w690162;

	wire w720162;

	wire w940162;

	wire w970162;

	wire w990162;

	wire w1020162;

	wire w1060162;

	wire w590163;

	wire w610163;

	wire w630163;

	wire w650163;

	wire w680163;

	wire w710163;

	wire w730163;

	wire w930163;

	wire w950163;

	wire w980163;

	wire w1010163;

	wire w1030163;

	wire w1050163;

	wire w1070163;

	wire w640164;

	wire w1020164;

	wire w600165;

	wire w640165;

	wire w650165;

	wire w690165;

	wire w710165;

	wire w730165;

	wire w930165;

	wire w950165;

	wire w970165;

	wire w1010165;

	wire w1020165;

	wire w1060165;

	wire w550167;
	repeater #(1, 1'b1, 0, 0) c550167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550167));
	wire w600167;
	repeater #(1, 1'b1, 0, 0) c600167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600167));
	wire w650167;
	repeater #(1, 1'b1, 0, 0) c650167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650167));
	wire w1010167;
	repeater #(1, 1'b0, 0, 0) c1010167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010167));
	wire w1060167;
	repeater #(1, 1'b1, 0, 0) c1060167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060167));
	wire w1110167;
	repeater #(1, 1'b1, 0, 0) c1110167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110167));
	wire w540168;

	wire w550168;
	repeater #(1, 1'b1, 0, 0) c550168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550168));
	wire w590168;

	wire w600168;
	repeater #(1, 1'b1, 0, 0) c600168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600168));
	wire w640168;

	wire w650168;
	repeater #(1, 1'b1, 0, 0) c650168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650168));
	wire w1010168;
	repeater #(1, 1'b0, 0, 0) c1010168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010168));
	wire w1020168;

	wire w1060168;
	repeater #(1, 1'b1, 0, 0) c1060168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060168));
	wire w1070168;

	wire w1110168;
	repeater #(1, 1'b1, 0, 0) c1110168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110168));
	wire w1120168;

	wire w1980169;

	wire w240170;

	wire w1960170;
	repeater #(1, 1'b1, 0, 0) c1960170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1960170));
	wire w40171;
	repeater #(1, 1'b1, 0, 0) c40171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40171));
	wire w220171;
	repeater #(1, 1'b1, 0, 0) c220171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220171));
	wire w380171;
	repeater #(1, 1'b1, 0, 0) c380171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380171));
	wire w550171;
	repeater #(1, 1'b1, 0, 0) c550171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550171));
	wire w600171;
	repeater #(1, 1'b1, 0, 0) c600171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600171));
	wire w650171;
	repeater #(1, 1'b0, 0, 0) c650171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650171));
	wire w1010171;
	repeater #(1, 1'b0, 0, 0) c1010171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010171));
	wire w1060171;
	repeater #(1, 1'b1, 0, 0) c1060171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060171));
	wire w1110171;
	repeater #(1, 1'b1, 0, 0) c1110171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110171));
	wire w1870171;
	repeater #(1, 1'b1, 0, 0) c1870171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870171));
	wire w2030171;
	repeater #(1, 1'b1, 0, 0) c2030171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030171));
	wire w130172;
	repeater #(1, 1'b1, 0, 0) c130172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130172));
	wire w290172;
	repeater #(1, 1'b1, 0, 0) c290172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290172));
	wire w540172;

	wire w550172;
	repeater #(1, 1'b1, 0, 0) c550172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550172));
	wire w590172;

	wire w600172;
	repeater #(1, 1'b0, 0, 0) c600172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600172));
	wire w640172;

	wire w650172;
	repeater #(1, 1'b0, 0, 0) c650172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650172));
	wire w1010172;
	repeater #(1, 1'b0, 0, 0) c1010172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010172));
	wire w1020172;

	wire w1060172;
	repeater #(1, 1'b1, 0, 0) c1060172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060172));
	wire w1070172;

	wire w1110172;
	repeater #(1, 1'b1, 0, 0) c1110172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110172));
	wire w1120172;

	wire w1240172;
	repeater #(1, 1'b0, 0, 0) c1240172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240172));
	wire w1440172;
	repeater #(1, 1'b0, 0, 0) c1440172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1440172));
	wire w1980172;

	wire w60173;

	wire w240173;

	wire w400173;

	wire w1900173;

	wire w2060173;

	wire w160174;

	wire w320174;

	wire w1870174;

	wire w1930174;

	wire w2010174;

	wire w2030174;

	wire w2040174;

	wire w10175;

	wire w90175;

	wire w130175;

	wire w190175;

	wire w270175;

	wire w290175;

	wire w300175;

	wire w350175;

	wire w430175;

	wire w550175;
	repeater #(1, 1'b0, 0, 0) c550175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550175));
	wire w600175;
	repeater #(1, 1'b0, 0, 0) c600175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600175));
	wire w650175;
	repeater #(1, 1'b0, 0, 0) c650175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650175));
	wire w1010175;
	repeater #(1, 1'b0, 0, 0) c1010175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010175));
	wire w1060175;
	repeater #(1, 1'b1, 0, 0) c1060175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060175));
	wire w1110175;
	repeater #(1, 1'b1, 0, 0) c1110175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110175));
	wire w60176;

	wire w400176;

	wire w540176;

	wire w550176;
	repeater #(1, 1'b0, 0, 0) c550176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550176));
	wire w590176;

	wire w600176;
	repeater #(1, 1'b0, 0, 0) c600176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600176));
	wire w640176;

	wire w650176;
	repeater #(1, 1'b0, 0, 0) c650176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650176));
	wire w1010176;
	repeater #(1, 1'b0, 0, 0) c1010176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010176));
	wire w1020176;

	wire w1060176;
	repeater #(1, 1'b1, 0, 0) c1060176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060176));
	wire w1070176;

	wire w1110176;
	repeater #(1, 1'b1, 0, 0) c1110176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110176));
	wire w1120176;

	wire w1950176;

	wire w1960176;

	wire w30177;

	wire w40177;

	wire w210177;

	wire w220177;

	wire w370177;

	wire w380177;

	wire w1870178;

	wire w1880178;

	wire w2010178;

	wire w2030178;

	wire w2040178;

	wire w910;

	wire w1310;

	wire w1410;

	wire w2710;

	wire w2910;

	wire w3010;

	wire w4310;

	wire w5510;
	repeater #(1, 1'b0, 0, 0) c5510 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5510));
	wire w6010;
	repeater #(1, 1'b0, 0, 0) c6010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6010));
	wire w6510;
	repeater #(1, 1'b0, 0, 0) c6510 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6510));
	wire w8110;

	wire w10110;
	repeater #(1, 1'b0, 0, 0) c10110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10110));
	wire w10610;
	repeater #(1, 1'b1, 0, 0) c10610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10610));
	wire w11110;
	repeater #(1, 1'b1, 0, 0) c11110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11110));
	wire w5411;

	wire w5511;
	repeater #(1, 1'b0, 0, 0) c5511 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5511));
	wire w5911;

	wire w6011;
	repeater #(1, 1'b0, 0, 0) c6011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6011));
	wire w6411;

	wire w6511;
	repeater #(1, 1'b0, 0, 0) c6511 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6511));
	wire w7211;
	repeater #(1, 1'b0, 0, 0) c7211 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7211));
	wire w9411;
	repeater #(1, 1'b0, 0, 0) c9411 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9411));
	wire w10111;
	repeater #(1, 1'b0, 0, 0) c10111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10111));
	wire w10211;

	wire w10611;
	repeater #(1, 1'b0, 0, 0) c10611 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10611));
	wire w10711;

	wire w11111;
	repeater #(1, 1'b0, 0, 0) c11111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11111));
	wire w11211;

	wire w19811;
	torch #(1'b1) c19811 (.i_clk(tick), .i_in(), .o_out(w19811));
	wire w19911;

	wire w612;
	torch #(1'b1) c612 (.i_clk(tick), .i_in(), .o_out(w612));
	wire w712;

	wire w2412;
	torch #(1'b1) c2412 (.i_clk(tick), .i_in(), .o_out(w2412));
	wire w2512;

	wire w4012;
	torch #(1'b1) c4012 (.i_clk(tick), .i_in(), .o_out(w4012));
	wire w4112;

	wire w6512;
	repeater #(2, 1'b0, 0, 0) c6512 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6512));
	wire w10112;
	repeater #(2, 1'b0, 0, 0) c10112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10112));
	wire w19912;

	wire w20112;

	wire w713;

	wire w913;

	wire w2513;

	wire w2713;

	wire w4113;

	wire w4313;

	wire w5413;

	wire w5513;

	wire w8313;
	assign w8313 = inputs[12];
	wire w11113;

	wire w11213;

	wire w5814;
	repeater #(2, 1'b0, 0, 0) c5814 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5814));
	wire w5914;
	repeater #(2, 1'b0, 0, 0) c5914 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5914));
	wire w6114;

	wire w10514;

	wire w10714;
	repeater #(2, 1'b0, 0, 0) c10714 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10714));
	wire w10814;
	repeater #(2, 1'b0, 0, 0) c10814 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10814));
	wire w20114;

	wire w20214;

	wire w20314;

	wire w915;

	wire w1015;

	wire w1115;

	wire w2715;

	wire w2815;

	wire w2915;

	wire w4315;

	wire w4415;

	wire w4515;

	wire w5915;

	wire w6115;
	repeater #(1, 1'b1, 0, 0) c6115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6115));
	wire w10515;
	repeater #(1, 1'b1, 0, 0) c10515 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10515));
	wire w10715;

	wire w19615;

	wire w19715;

	wire w20315;

	wire w416;

	wire w516;

	wire w1116;

	wire w2216;

	wire w2316;

	wire w2916;

	wire w3816;

	wire w3916;

	wire w4516;

	wire w5516;

	wire w5916;

	wire w10716;

	wire w11116;

	wire w5517;

	wire w5717;
	repeater #(1, 1'b1, 0, 0) c5717 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5717));
	wire w6217;

	wire w6617;

	wire w10017;

	wire w10417;

	wire w10917;
	repeater #(1, 1'b0, 0, 0) c10917 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10917));
	wire w11117;

	wire w19317;
	torch #(1'b0) c19317 (.i_clk(tick), .i_in(), .o_out(w19317));
	wire w20117;
	repeater #(1, 1'b0, 0, 0) c20117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20117));
	wire w20317;
	torch #(1'b0) c20317 (.i_clk(tick), .i_in(), .o_out(w20317));
	wire w118;
	torch #(1'b0) c118 (.i_clk(tick), .i_in(), .o_out(w118));
	wire w918;
	repeater #(1, 1'b0, 0, 0) c918 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w918));
	wire w1118;
	torch #(1'b0) c1118 (.i_clk(tick), .i_in(), .o_out(w1118));
	wire w1918;
	torch #(1'b0) c1918 (.i_clk(tick), .i_in(), .o_out(w1918));
	wire w2718;
	repeater #(1, 1'b0, 0, 0) c2718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2718));
	wire w2918;
	torch #(1'b0) c2918 (.i_clk(tick), .i_in(), .o_out(w2918));
	wire w3518;
	torch #(1'b0) c3518 (.i_clk(tick), .i_in(), .o_out(w3518));
	wire w4318;
	repeater #(1, 1'b0, 0, 0) c4318 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4318));
	wire w4518;
	torch #(1'b0) c4518 (.i_clk(tick), .i_in(), .o_out(w4518));
	wire w6218;

	wire w6418;
	repeater #(1, 1'b0, 0, 0) c6418 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6418));
	wire w6518;

	wire w10118;

	wire w10218;
	repeater #(1, 1'b1, 0, 0) c10218 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10218));
	wire w10418;

	wire w5819;

	wire w10819;

	wire w12419;
	repeater #(1, 1'b0, 0, 0) c12419 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12419));
	wire w14419;
	repeater #(1, 1'b0, 0, 0) c14419 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14419));
	wire w20519;
	repeater #(1, 1'b1, 0, 0) c20519 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20519));
	wire w31110;
	repeater #(1, 1'b1, 0, 0) c31110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31110));
	wire w55110;

	wire w56110;
	repeater #(1, 1'b0, 0, 0) c56110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56110));
	wire w63110;
	repeater #(2, 1'b1, 0, 0) c63110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63110));
	wire w103110;
	repeater #(2, 1'b1, 0, 0) c103110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103110));
	wire w110110;
	repeater #(1, 1'b1, 0, 0) c110110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110110));
	wire w111110;

	wire w202111;
	torch #(1'b1) c202111 (.i_clk(tick), .i_in(), .o_out(w202111));
	wire w10112;
	torch #(1'b1) c10112 (.i_clk(tick), .i_in(), .o_out(w10112));
	wire w28112;
	torch #(1'b1) c28112 (.i_clk(tick), .i_in(), .o_out(w28112));
	wire w44112;
	torch #(1'b1) c44112 (.i_clk(tick), .i_in(), .o_out(w44112));
	wire w194113;
	torch #(1'b1) c194113 (.i_clk(tick), .i_in(), .o_out(w194113));
	wire w2114;
	torch #(1'b1) c2114 (.i_clk(tick), .i_in(), .o_out(w2114));
	wire w20114;
	torch #(1'b1) c20114 (.i_clk(tick), .i_in(), .o_out(w20114));
	wire w36114;
	torch #(1'b1) c36114 (.i_clk(tick), .i_in(), .o_out(w36114));
	wire w201114;
	repeater #(1, 1'b0, 0, 0) c201114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201114));
	wire w9115;
	repeater #(1, 1'b0, 0, 0) c9115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9115));
	wire w27115;
	repeater #(1, 1'b0, 0, 0) c27115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27115));
	wire w43115;
	repeater #(1, 1'b0, 0, 0) c43115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43115));
	wire w195115;
	repeater #(1, 1'b0, 0, 0) c195115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195115));
	wire w3116;
	repeater #(1, 1'b0, 0, 0) c3116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3116));
	wire w21116;
	repeater #(1, 1'b0, 0, 0) c21116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21116));
	wire w37116;
	repeater #(1, 1'b0, 0, 0) c37116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37116));
	wire w124125;
	repeater #(1, 1'b0, 0, 0) c124125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124125));
	wire w144125;
	repeater #(1, 1'b0, 0, 0) c144125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144125));
	wire w124141;
	repeater #(1, 1'b0, 0, 0) c124141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124141));
	wire w144141;
	repeater #(1, 1'b0, 0, 0) c144141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144141));
	wire w121162;
	torch #(1'b1) c121162 (.i_clk(tick), .i_in(), .o_out(w121162));
	wire w125162;
	torch #(1'b1) c125162 (.i_clk(tick), .i_in(), .o_out(w125162));
	wire w129162;
	torch #(1'b0) c129162 (.i_clk(tick), .i_in(), .o_out(w129162));
	wire w133162;
	torch #(1'b1) c133162 (.i_clk(tick), .i_in(), .o_out(w133162));
	wire w137162;
	torch #(1'b0) c137162 (.i_clk(tick), .i_in(), .o_out(w137162));
	wire w141162;
	torch #(1'b1) c141162 (.i_clk(tick), .i_in(), .o_out(w141162));
	wire w145162;
	torch #(1'b1) c145162 (.i_clk(tick), .i_in(), .o_out(w145162));
	wire w119163;
	torch #(1'b1) c119163 (.i_clk(tick), .i_in(), .o_out(w119163));
	wire w123163;
	torch #(1'b1) c123163 (.i_clk(tick), .i_in(), .o_out(w123163));
	wire w127163;
	torch #(1'b1) c127163 (.i_clk(tick), .i_in(), .o_out(w127163));
	wire w131163;
	torch #(1'b1) c131163 (.i_clk(tick), .i_in(), .o_out(w131163));
	wire w135163;
	torch #(1'b1) c135163 (.i_clk(tick), .i_in(), .o_out(w135163));
	wire w139163;
	torch #(1'b1) c139163 (.i_clk(tick), .i_in(), .o_out(w139163));
	wire w143163;
	torch #(1'b1) c143163 (.i_clk(tick), .i_in(), .o_out(w143163));
	wire w121166;
	torch #(1'b1) c121166 (.i_clk(tick), .i_in(), .o_out(w121166));
	wire w125166;
	torch #(1'b1) c125166 (.i_clk(tick), .i_in(), .o_out(w125166));
	wire w129166;
	torch #(1'b1) c129166 (.i_clk(tick), .i_in(), .o_out(w129166));
	wire w133166;
	torch #(1'b0) c133166 (.i_clk(tick), .i_in(), .o_out(w133166));
	wire w137166;
	torch #(1'b1) c137166 (.i_clk(tick), .i_in(), .o_out(w137166));
	wire w141166;
	torch #(1'b1) c141166 (.i_clk(tick), .i_in(), .o_out(w141166));
	wire w145166;
	torch #(1'b1) c145166 (.i_clk(tick), .i_in(), .o_out(w145166));
	wire w120174;
	torch #(1'b1) c120174 (.i_clk(tick), .i_in(), .o_out(w120174));
	wire w124174;
	torch #(1'b1) c124174 (.i_clk(tick), .i_in(), .o_out(w124174));
	wire w128174;
	torch #(1'b1) c128174 (.i_clk(tick), .i_in(), .o_out(w128174));
	wire w132174;
	torch #(1'b1) c132174 (.i_clk(tick), .i_in(), .o_out(w132174));
	wire w136174;
	torch #(1'b1) c136174 (.i_clk(tick), .i_in(), .o_out(w136174));
	wire w140174;
	torch #(1'b1) c140174 (.i_clk(tick), .i_in(), .o_out(w140174));
	wire w144174;
	torch #(1'b1) c144174 (.i_clk(tick), .i_in(), .o_out(w144174));
	wire w154176;
	repeater #(1, 1'b0, 0, 0) c154176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154176));
	wire w1211107;
	repeater #(1, 1'b0, 0, 0) c1211107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1211107));
	wire w1251107;
	repeater #(1, 1'b0, 0, 0) c1251107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1251107));
	wire w1291107;
	repeater #(1, 1'b0, 0, 0) c1291107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1291107));
	wire w1331107;
	repeater #(1, 1'b1, 0, 0) c1331107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1331107));
	wire w1371107;
	repeater #(1, 1'b0, 0, 0) c1371107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1371107));
	wire w1411107;
	repeater #(1, 1'b0, 0, 0) c1411107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1411107));
	wire w1451107;
	repeater #(1, 1'b0, 0, 0) c1451107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1451107));
	wire w1211110;
	torch #(1'b1) c1211110 (.i_clk(tick), .i_in(), .o_out(w1211110));
	wire w1251110;
	torch #(1'b1) c1251110 (.i_clk(tick), .i_in(), .o_out(w1251110));
	wire w1291110;
	torch #(1'b1) c1291110 (.i_clk(tick), .i_in(), .o_out(w1291110));
	wire w1331110;
	torch #(1'b0) c1331110 (.i_clk(tick), .i_in(), .o_out(w1331110));
	wire w1371110;
	torch #(1'b1) c1371110 (.i_clk(tick), .i_in(), .o_out(w1371110));
	wire w1411110;
	torch #(1'b1) c1411110 (.i_clk(tick), .i_in(), .o_out(w1411110));
	wire w1451110;
	torch #(1'b1) c1451110 (.i_clk(tick), .i_in(), .o_out(w1451110));
	wire w1321113;
	repeater #(1, 1'b0, 0, 0) c1321113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321113));
	wire w1341113;
	repeater #(1, 1'b0, 0, 0) c1341113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1341113));
	wire w1361113;
	repeater #(1, 1'b1, 0, 0) c1361113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361113));
	wire w1381113;
	repeater #(1, 1'b1, 0, 0) c1381113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1381113));
	wire w1401113;
	repeater #(1, 1'b1, 0, 0) c1401113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401113));
	wire w1421113;
	repeater #(1, 1'b1, 0, 0) c1421113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1421113));
	wire w1441113;
	repeater #(1, 1'b1, 0, 0) c1441113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441113));
	wire w1461113;
	repeater #(1, 1'b1, 0, 0) c1461113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1461113));
	wire w1301115;
	repeater #(1, 1'b1, 0, 0) c1301115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1301115));
	wire w1281117;
	repeater #(1, 1'b1, 0, 0) c1281117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281117));
	wire w1261119;
	repeater #(1, 1'b1, 0, 0) c1261119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1261119));
	wire w1241121;
	repeater #(1, 1'b1, 0, 0) c1241121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241121));
	wire w1221123;
	repeater #(1, 1'b1, 0, 0) c1221123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221123));
	wire w1201125;
	repeater #(1, 1'b1, 0, 0) c1201125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201125));
	wire w101131;
	torch #(1'b1) c101131 (.i_clk(tick), .i_in(), .o_out(w101131));
	wire w441131;
	repeater #(1, 1'b1, 0, 0) c441131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w441131));
	wire w781131;
	torch #(1'b1) c781131 (.i_clk(tick), .i_in(), .o_out(w781131));
	wire w1121131;
	repeater #(1, 1'b1, 0, 0) c1121131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121131));
	wire w81133;
	repeater #(1, 1'b1, 0, 0) c81133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81133));
	wire w421133;
	repeater #(1, 1'b1, 0, 0) c421133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w421133));
	wire w761133;
	repeater #(1, 1'b1, 0, 0) c761133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w761133));
	wire w1101133;
	repeater #(1, 1'b1, 0, 0) c1101133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101133));
	wire w1461134;
	repeater #(1, 1'b1, 0, 0) c1461134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1461134));
	wire w61135;
	torch #(1'b1) c61135 (.i_clk(tick), .i_in(), .o_out(w61135));
	wire w401135;
	repeater #(1, 1'b1, 0, 0) c401135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w401135));
	wire w741135;
	torch #(1'b1) c741135 (.i_clk(tick), .i_in(), .o_out(w741135));
	wire w1081135;
	repeater #(1, 1'b1, 0, 0) c1081135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081135));
	wire w12800;
	repeater #(1, 1'b1, 0, 0) c12800 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12800));
	wire w19600;
	repeater #(1, 1'b1, 0, 0) c19600 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19600));
	wire w2201;
	repeater #(1, 1'b1, 0, 0) c2201 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2201));
	wire w5601;
	repeater #(1, 1'b1, 0, 0) c5601 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5601));
	wire w9001;
	repeater #(1, 1'b1, 0, 0) c9001 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9001));
	wire w12602;
	repeater #(1, 1'b1, 0, 0) c12602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12602));
	wire w19402;
	torch #(1'b1) c19402 (.i_clk(tick), .i_in(), .o_out(w19402));
	wire w2003;
	repeater #(1, 1'b1, 0, 0) c2003 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2003));
	wire w5403;
	torch #(1'b1) c5403 (.i_clk(tick), .i_in(), .o_out(w5403));
	wire w8803;
	repeater #(1, 1'b1, 0, 0) c8803 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8803));
	wire w12404;
	repeater #(1, 1'b1, 0, 0) c12404 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12404));
	wire w19204;
	repeater #(1, 1'b1, 0, 0) c19204 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19204));
	wire w1805;
	repeater #(1, 1'b1, 0, 0) c1805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1805));
	wire w5205;
	repeater #(1, 1'b1, 0, 0) c5205 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5205));
	wire w8605;
	repeater #(1, 1'b1, 0, 0) c8605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8605));
	wire w17605;
	repeater #(1, 1'b1, 0, 0) c17605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17605));
	wire w17805;
	torch #(1'b1) c17805 (.i_clk(tick), .i_in(), .o_out(w17805));
	wire w18005;
	repeater #(1, 1'b1, 0, 0) c18005 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18005));
	wire w18205;
	torch #(1'b1) c18205 (.i_clk(tick), .i_in(), .o_out(w18205));
	wire w18405;
	repeater #(1, 1'b1, 0, 0) c18405 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18405));
	wire w18605;
	torch #(1'b1) c18605 (.i_clk(tick), .i_in(), .o_out(w18605));
	wire w18805;
	repeater #(1, 1'b0, 0, 0) c18805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18805));
	wire w19005;
	torch #(1'b0) c19005 (.i_clk(tick), .i_in(), .o_out(w19005));
	wire w206;
	repeater #(1, 1'b1, 0, 0) c206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206));
	wire w406;
	repeater #(1, 1'b1, 0, 0) c406 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w406));
	wire w606;
	repeater #(1, 1'b1, 0, 0) c606 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w606));
	wire w806;
	repeater #(1, 1'b1, 0, 0) c806 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w806));
	wire w1006;
	repeater #(1, 1'b1, 0, 0) c1006 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1006));
	wire w1206;
	repeater #(1, 1'b1, 0, 0) c1206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1206));
	wire w1406;
	repeater #(1, 1'b0, 0, 0) c1406 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1406));
	wire w1606;
	repeater #(1, 1'b0, 0, 0) c1606 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1606));
	wire w3806;
	torch #(1'b1) c3806 (.i_clk(tick), .i_in(), .o_out(w3806));
	wire w4206;
	torch #(1'b1) c4206 (.i_clk(tick), .i_in(), .o_out(w4206));
	wire w4606;
	torch #(1'b1) c4606 (.i_clk(tick), .i_in(), .o_out(w4606));
	wire w5006;
	torch #(1'b0) c5006 (.i_clk(tick), .i_in(), .o_out(w5006));
	wire w7006;
	repeater #(1, 1'b1, 0, 0) c7006 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7006));
	wire w7206;
	repeater #(1, 1'b1, 0, 0) c7206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7206));
	wire w7406;
	repeater #(1, 1'b1, 0, 0) c7406 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7406));
	wire w7606;
	repeater #(1, 1'b1, 0, 0) c7606 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7606));
	wire w7806;
	repeater #(1, 1'b1, 0, 0) c7806 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7806));
	wire w8006;
	repeater #(1, 1'b1, 0, 0) c8006 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8006));
	wire w8206;
	repeater #(1, 1'b0, 0, 0) c8206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8206));
	wire w8406;
	repeater #(1, 1'b0, 0, 0) c8406 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8406));
	wire w12206;
	repeater #(1, 1'b1, 0, 0) c12206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12206));
	wire w3707;
	repeater #(1, 1'b1, 0, 0) c3707 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3707));
	wire w4107;
	repeater #(1, 1'b1, 0, 0) c4107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4107));
	wire w4507;
	repeater #(1, 1'b1, 0, 0) c4507 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4507));
	wire w4907;
	repeater #(1, 1'b0, 0, 0) c4907 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4907));
	wire w10807;
	repeater #(1, 1'b1, 0, 0) c10807 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10807));
	wire w11007;
	repeater #(1, 1'b1, 0, 0) c11007 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11007));
	wire w11207;
	repeater #(1, 1'b1, 0, 0) c11207 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11207));
	wire w11407;
	repeater #(1, 1'b1, 0, 0) c11407 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11407));
	wire w11607;
	repeater #(1, 1'b0, 0, 0) c11607 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11607));
	wire w11807;
	repeater #(1, 1'b0, 0, 0) c11807 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11807));
	wire w12007;
	repeater #(1, 1'b1, 0, 0) c12007 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12007));
	wire w3809;
	torch #(1'b1) c3809 (.i_clk(tick), .i_in(), .o_out(w3809));
	wire w4209;
	torch #(1'b1) c4209 (.i_clk(tick), .i_in(), .o_out(w4209));
	wire w4609;
	torch #(1'b1) c4609 (.i_clk(tick), .i_in(), .o_out(w4609));
	wire w5009;
	torch #(1'b1) c5009 (.i_clk(tick), .i_in(), .o_out(w5009));
	wire w5409;
	torch #(1'b1) c5409 (.i_clk(tick), .i_in(), .o_out(w5409));
	wire w5809;
	torch #(1'b1) c5809 (.i_clk(tick), .i_in(), .o_out(w5809));
	wire w6209;
	torch #(1'b1) c6209 (.i_clk(tick), .i_in(), .o_out(w6209));
	wire w7209;
	torch #(1'b1) c7209 (.i_clk(tick), .i_in(), .o_out(w7209));
	wire w7609;
	torch #(1'b1) c7609 (.i_clk(tick), .i_in(), .o_out(w7609));
	wire w8009;
	torch #(1'b1) c8009 (.i_clk(tick), .i_in(), .o_out(w8009));
	wire w8409;
	torch #(1'b0) c8409 (.i_clk(tick), .i_in(), .o_out(w8409));
	wire w8809;
	torch #(1'b1) c8809 (.i_clk(tick), .i_in(), .o_out(w8809));
	wire w9209;
	torch #(1'b1) c9209 (.i_clk(tick), .i_in(), .o_out(w9209));
	wire w9609;
	torch #(1'b1) c9609 (.i_clk(tick), .i_in(), .o_out(w9609));
	wire w17609;
	repeater #(2, 1'b1, 0, 0) c17609 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17609));
	wire w18009;
	repeater #(2, 1'b1, 0, 0) c18009 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18009));
	wire w18409;
	repeater #(2, 1'b1, 0, 0) c18409 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18409));
	wire w20009;
	repeater #(2, 1'b1, 0, 0) c20009 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20009));
	wire w2010;
	repeater #(2, 1'b1, 0, 0) c2010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010));
	wire w6010;
	repeater #(2, 1'b1, 0, 0) c6010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6010));
	wire w10010;
	repeater #(2, 1'b1, 0, 0) c10010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10010));
	wire w26010;
	repeater #(2, 1'b1, 0, 0) c26010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26010));
	wire w43011;
	torch #(1'b0) c43011 (.i_clk(tick), .i_in(), .o_out(w43011));
	wire w47011;
	torch #(1'b0) c47011 (.i_clk(tick), .i_in(), .o_out(w47011));
	wire w51011;
	torch #(1'b0) c51011 (.i_clk(tick), .i_in(), .o_out(w51011));
	wire w55011;
	torch #(1'b0) c55011 (.i_clk(tick), .i_in(), .o_out(w55011));
	wire w79011;
	torch #(1'b1) c79011 (.i_clk(tick), .i_in(), .o_out(w79011));
	wire w83011;
	torch #(1'b1) c83011 (.i_clk(tick), .i_in(), .o_out(w83011));
	wire w87011;
	torch #(1'b1) c87011 (.i_clk(tick), .i_in(), .o_out(w87011));
	wire w91011;
	torch #(1'b1) c91011 (.i_clk(tick), .i_in(), .o_out(w91011));
	wire w176011;
	torch #(1'b1) c176011 (.i_clk(tick), .i_in(), .o_out(w176011));
	wire w186011;
	repeater #(1, 1'b1, 0, 0) c186011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186011));
	wire w192011;
	torch #(1'b1) c192011 (.i_clk(tick), .i_in(), .o_out(w192011));
	wire w202011;
	repeater #(1, 1'b1, 0, 0) c202011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202011));
	wire w2012;
	torch #(1'b1) c2012 (.i_clk(tick), .i_in(), .o_out(w2012));
	wire w12012;
	repeater #(1, 1'b1, 0, 0) c12012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12012));
	wire w18012;
	torch #(1'b1) c18012 (.i_clk(tick), .i_in(), .o_out(w18012));
	wire w28012;
	repeater #(1, 1'b1, 0, 0) c28012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28012));
	wire w177014;
	repeater #(1, 1'b1, 0, 0) c177014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177014));
	wire w193014;
	repeater #(1, 1'b1, 0, 0) c193014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193014));
	wire w3015;
	repeater #(1, 1'b1, 0, 0) c3015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3015));
	wire w19015;
	repeater #(1, 1'b1, 0, 0) c19015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19015));
	wire w186015;
	repeater #(1, 1'b1, 0, 0) c186015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186015));
	wire w202015;
	repeater #(1, 1'b1, 0, 0) c202015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202015));
	wire w12016;
	repeater #(1, 1'b1, 0, 0) c12016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12016));
	wire w28016;
	repeater #(1, 1'b1, 0, 0) c28016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28016));
	wire w175016;

	wire w191016;

	wire w1017;

	wire w17017;

	wire w106017;
	repeater #(1, 1'b1, 0, 0) c106017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106017));
	wire w110017;
	repeater #(1, 1'b1, 0, 0) c110017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110017));
	wire w114017;
	repeater #(1, 1'b1, 0, 0) c114017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114017));
	wire w118017;
	repeater #(1, 1'b1, 0, 0) c118017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118017));
	wire w122017;
	repeater #(1, 1'b1, 0, 0) c122017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122017));
	wire w126017;
	repeater #(1, 1'b1, 0, 0) c126017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126017));
	wire w130017;
	repeater #(1, 1'b1, 0, 0) c130017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130017));
	wire w183017;

	wire w199017;

	wire w9018;

	wire w25018;

	wire w180018;

	wire w185018;

	wire w186018;

	wire w196018;

	wire w202018;

	wire w6019;

	wire w11019;

	wire w12019;

	wire w22019;

	wire w28019;

	wire w175019;

	wire w1020;

	wire w178020;

	wire w194020;

	wire w4021;

	wire w20021;

	wire w133021;
	repeater #(1, 1'b0, 0, 0) c133021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133021));
	wire w184021;

	wire w185021;

	wire w200021;

	wire w201021;

	wire w10022;

	wire w11022;

	wire w26022;

	wire w27022;

	wire w194022;

	wire w198022;

	wire w20023;

	wire w24023;

	wire w103023;
	repeater #(1, 1'b0, 0, 0) c103023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103023));
	wire w112026;
	torch #(1'b1) c112026 (.i_clk(tick), .i_in(), .o_out(w112026));
	wire w116026;
	torch #(1'b1) c116026 (.i_clk(tick), .i_in(), .o_out(w116026));
	wire w120026;
	torch #(1'b1) c120026 (.i_clk(tick), .i_in(), .o_out(w120026));
	wire w124026;
	torch #(1'b1) c124026 (.i_clk(tick), .i_in(), .o_out(w124026));
	wire w175026;

	wire w176026;

	wire w179026;

	wire w180026;

	wire w183026;

	wire w184026;

	wire w187026;

	wire w188026;

	wire w191026;

	wire w192026;

	wire w195026;

	wire w196026;

	wire w199026;

	wire w200026;

	wire w1027;

	wire w2027;

	wire w5027;

	wire w6027;

	wire w9027;

	wire w10027;

	wire w13027;

	wire w14027;

	wire w17027;

	wire w18027;

	wire w21027;

	wire w22027;

	wire w25027;

	wire w26027;

	wire w176028;

	wire w180028;

	wire w184028;

	wire w188028;

	wire w192028;

	wire w196028;

	wire w200028;

	wire w2029;

	wire w6029;

	wire w10029;

	wire w14029;

	wire w18029;

	wire w22029;

	wire w26029;

	wire w105030;
	torch #(1'b0) c105030 (.i_clk(tick), .i_in(), .o_out(w105030));
	wire w109030;
	torch #(1'b0) c109030 (.i_clk(tick), .i_in(), .o_out(w109030));
	wire w113030;
	torch #(1'b0) c113030 (.i_clk(tick), .i_in(), .o_out(w113030));
	wire w117030;
	torch #(1'b0) c117030 (.i_clk(tick), .i_in(), .o_out(w117030));
	wire w121030;
	torch #(1'b0) c121030 (.i_clk(tick), .i_in(), .o_out(w121030));
	wire w125030;
	torch #(1'b0) c125030 (.i_clk(tick), .i_in(), .o_out(w125030));
	wire w129030;
	torch #(1'b0) c129030 (.i_clk(tick), .i_in(), .o_out(w129030));
	wire w51031;

	wire w83031;

	wire w174031;

	wire w178031;

	wire w182031;

	wire w186031;

	wire w0032;

	wire w4032;

	wire w8032;

	wire w12032;

	wire w106032;
	torch #(1'b1) c106032 (.i_clk(tick), .i_in(), .o_out(w106032));
	wire w110032;
	torch #(1'b1) c110032 (.i_clk(tick), .i_in(), .o_out(w110032));
	wire w114032;
	torch #(1'b1) c114032 (.i_clk(tick), .i_in(), .o_out(w114032));
	wire w118032;
	torch #(1'b1) c118032 (.i_clk(tick), .i_in(), .o_out(w118032));
	wire w122032;
	torch #(1'b1) c122032 (.i_clk(tick), .i_in(), .o_out(w122032));
	wire w126032;
	torch #(1'b1) c126032 (.i_clk(tick), .i_in(), .o_out(w126032));
	wire w130032;
	torch #(1'b1) c130032 (.i_clk(tick), .i_in(), .o_out(w130032));
	wire w186033;

	wire w12034;

	wire w38034;

	wire w39034;
	repeater #(1, 1'b1, 0, 0) c39034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39034));
	wire w43034;

	wire w44034;
	repeater #(1, 1'b1, 0, 0) c44034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44034));
	wire w48034;

	wire w49034;
	repeater #(1, 1'b1, 0, 0) c49034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49034));
	wire w85034;
	repeater #(1, 1'b0, 0, 0) c85034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85034));
	wire w86034;

	wire w90034;
	repeater #(1, 1'b1, 0, 0) c90034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90034));
	wire w91034;

	wire w95034;
	repeater #(1, 1'b1, 0, 0) c95034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95034));
	wire w96034;

	wire w107034;
	torch #(1'b0) c107034 (.i_clk(tick), .i_in(), .o_out(w107034));
	wire w111034;
	torch #(1'b0) c111034 (.i_clk(tick), .i_in(), .o_out(w111034));
	wire w115034;
	torch #(1'b0) c115034 (.i_clk(tick), .i_in(), .o_out(w115034));
	wire w119034;
	torch #(1'b0) c119034 (.i_clk(tick), .i_in(), .o_out(w119034));
	wire w123034;
	torch #(1'b0) c123034 (.i_clk(tick), .i_in(), .o_out(w123034));
	wire w127034;
	torch #(1'b0) c127034 (.i_clk(tick), .i_in(), .o_out(w127034));
	wire w131034;
	torch #(1'b0) c131034 (.i_clk(tick), .i_in(), .o_out(w131034));
	wire w184034;
	repeater #(1, 1'b0, 0, 0) c184034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184034));
	wire w10035;
	repeater #(1, 1'b1, 0, 0) c10035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10035));
	wire w175035;
	repeater #(1, 1'b1, 0, 0) c175035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175035));
	wire w191035;
	repeater #(1, 1'b1, 0, 0) c191035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191035));
	wire w1036;
	repeater #(1, 1'b1, 0, 0) c1036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1036));
	wire w17036;
	repeater #(1, 1'b1, 0, 0) c17036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17036));
	wire w186036;

	wire w12037;

	wire w133037;
	repeater #(1, 1'b0, 0, 0) c133037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133037));
	wire w178037;

	wire w194037;

	wire w4038;

	wire w20038;

	wire w38038;

	wire w39038;
	repeater #(1, 1'b0, 0, 0) c39038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39038));
	wire w43038;

	wire w44038;
	repeater #(1, 1'b0, 0, 0) c44038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44038));
	wire w48038;

	wire w49038;
	repeater #(1, 1'b0, 0, 0) c49038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49038));
	wire w85038;
	repeater #(1, 1'b0, 0, 0) c85038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85038));
	wire w86038;

	wire w90038;
	repeater #(1, 1'b1, 0, 0) c90038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90038));
	wire w91038;

	wire w95038;
	repeater #(1, 1'b1, 0, 0) c95038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95038));
	wire w96038;

	wire w175038;

	wire w176038;

	wire w181038;

	wire w189038;

	wire w191038;

	wire w192038;

	wire w197038;

	wire w1039;

	wire w2039;

	wire w7039;

	wire w15039;

	wire w17039;

	wire w18039;

	wire w23039;

	wire w103039;
	repeater #(1, 1'b0, 0, 0) c103039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103039));
	wire w183040;

	wire w184040;

	wire w199040;

	wire w200040;

	wire w9041;

	wire w10041;

	wire w25041;

	wire w26041;

	wire w38042;

	wire w39042;
	repeater #(1, 1'b0, 0, 0) c39042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39042));
	wire w43042;

	wire w44042;
	repeater #(1, 1'b0, 0, 0) c44042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44042));
	wire w48042;

	wire w49042;
	repeater #(1, 1'b0, 0, 0) c49042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49042));
	wire w85042;
	repeater #(1, 1'b0, 0, 0) c85042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85042));
	wire w86042;

	wire w90042;
	repeater #(1, 1'b1, 0, 0) c90042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90042));
	wire w91042;

	wire w95042;
	repeater #(1, 1'b1, 0, 0) c95042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95042));
	wire w96042;

	wire w112042;
	torch #(1'b1) c112042 (.i_clk(tick), .i_in(), .o_out(w112042));
	wire w116042;
	torch #(1'b1) c116042 (.i_clk(tick), .i_in(), .o_out(w116042));
	wire w120042;
	torch #(1'b1) c120042 (.i_clk(tick), .i_in(), .o_out(w120042));
	wire w124042;
	torch #(1'b1) c124042 (.i_clk(tick), .i_in(), .o_out(w124042));
	wire w175042;

	wire w176042;

	wire w189042;

	wire w191042;

	wire w192042;

	wire w1043;

	wire w2043;

	wire w15043;

	wire w17043;

	wire w18043;

	wire w65044;
	repeater #(1, 1'b1, 0, 0) c65044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65044));
	wire w186044;
	torch #(1'b1) c186044 (.i_clk(tick), .i_in(), .o_out(w186044));
	wire w187044;

	wire w12045;
	torch #(1'b1) c12045 (.i_clk(tick), .i_in(), .o_out(w12045));
	wire w13045;

	wire w40045;
	repeater #(2, 1'b0, 0, 0) c40045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40045));
	wire w94045;
	repeater #(2, 1'b0, 0, 0) c94045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94045));
	wire w187045;

	wire w189045;

	wire w13046;

	wire w15046;

	wire w37046;
	repeater #(1, 1'b1, 0, 0) c37046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37046));
	wire w45046;
	repeater #(1, 1'b0, 0, 0) c45046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45046));
	wire w46046;
	repeater #(2, 1'b0, 0, 0) c46046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46046));
	wire w88046;
	repeater #(2, 1'b0, 0, 0) c88046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88046));
	wire w89046;
	repeater #(1, 1'b0, 0, 0) c89046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89046));
	wire w97046;
	repeater #(1, 1'b0, 0, 0) c97046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97046));
	wire w105046;
	torch #(1'b0) c105046 (.i_clk(tick), .i_in(), .o_out(w105046));
	wire w109046;
	torch #(1'b0) c109046 (.i_clk(tick), .i_in(), .o_out(w109046));
	wire w113046;
	torch #(1'b0) c113046 (.i_clk(tick), .i_in(), .o_out(w113046));
	wire w117046;
	torch #(1'b1) c117046 (.i_clk(tick), .i_in(), .o_out(w117046));
	wire w121046;
	torch #(1'b0) c121046 (.i_clk(tick), .i_in(), .o_out(w121046));
	wire w125046;
	torch #(1'b0) c125046 (.i_clk(tick), .i_in(), .o_out(w125046));
	wire w129046;
	torch #(1'b0) c129046 (.i_clk(tick), .i_in(), .o_out(w129046));
	wire w41047;
	repeater #(1, 1'b0, 0, 0) c41047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41047));
	wire w66047;

	wire w93047;
	repeater #(1, 1'b0, 0, 0) c93047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93047));
	wire w189047;

	wire w190047;

	wire w191047;

	wire w15048;

	wire w16048;

	wire w17048;

	wire w47048;

	wire w51048;
	repeater #(1, 1'b0, 0, 0) c51048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51048));
	wire w67048;
	repeater #(2, 1'b0, 0, 0) c67048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67048));
	wire w83048;
	repeater #(1, 1'b0, 0, 0) c83048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83048));
	wire w87048;

	wire w106048;
	torch #(1'b1) c106048 (.i_clk(tick), .i_in(), .o_out(w106048));
	wire w110048;
	torch #(1'b1) c110048 (.i_clk(tick), .i_in(), .o_out(w110048));
	wire w114048;
	torch #(1'b1) c114048 (.i_clk(tick), .i_in(), .o_out(w114048));
	wire w118048;
	torch #(1'b1) c118048 (.i_clk(tick), .i_in(), .o_out(w118048));
	wire w122048;
	torch #(1'b1) c122048 (.i_clk(tick), .i_in(), .o_out(w122048));
	wire w126048;
	torch #(1'b1) c126048 (.i_clk(tick), .i_in(), .o_out(w126048));
	wire w130048;
	torch #(1'b1) c130048 (.i_clk(tick), .i_in(), .o_out(w130048));
	wire w184048;

	wire w185048;

	wire w191048;

	wire w200048;

	wire w201048;

	wire w10049;

	wire w11049;

	wire w17049;

	wire w26049;

	wire w27049;

	wire w48049;

	wire w57049;
	repeater #(2, 1'b0, 0, 0) c57049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57049));
	wire w77049;
	repeater #(2, 1'b1, 0, 0) c77049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77049));
	wire w86049;

	wire w47050;
	repeater #(2, 1'b1, 0, 0) c47050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47050));
	wire w58050;

	wire w76050;

	wire w87050;
	repeater #(2, 1'b0, 0, 0) c87050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87050));
	wire w107050;
	torch #(1'b0) c107050 (.i_clk(tick), .i_in(), .o_out(w107050));
	wire w111050;
	torch #(1'b0) c111050 (.i_clk(tick), .i_in(), .o_out(w111050));
	wire w115050;
	torch #(1'b0) c115050 (.i_clk(tick), .i_in(), .o_out(w115050));
	wire w119050;
	torch #(1'b0) c119050 (.i_clk(tick), .i_in(), .o_out(w119050));
	wire w123050;
	torch #(1'b0) c123050 (.i_clk(tick), .i_in(), .o_out(w123050));
	wire w127050;
	torch #(1'b0) c127050 (.i_clk(tick), .i_in(), .o_out(w127050));
	wire w131050;
	torch #(1'b0) c131050 (.i_clk(tick), .i_in(), .o_out(w131050));
	wire w181050;
	torch #(1'b0) c181050 (.i_clk(tick), .i_in(), .o_out(w181050));
	wire w189050;
	repeater #(1, 1'b1, 0, 0) c189050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189050));
	wire w191050;
	torch #(1'b0) c191050 (.i_clk(tick), .i_in(), .o_out(w191050));
	wire w197050;
	torch #(1'b0) c197050 (.i_clk(tick), .i_in(), .o_out(w197050));
	wire w7051;
	torch #(1'b0) c7051 (.i_clk(tick), .i_in(), .o_out(w7051));
	wire w15051;
	repeater #(1, 1'b1, 0, 0) c15051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15051));
	wire w17051;
	torch #(1'b0) c17051 (.i_clk(tick), .i_in(), .o_out(w17051));
	wire w23051;
	torch #(1'b0) c23051 (.i_clk(tick), .i_in(), .o_out(w23051));
	wire w41051;

	wire w42051;

	wire w92051;

	wire w93051;

	wire w40052;

	wire w49052;

	wire w85052;

	wire w94052;

	wire w177052;
	repeater #(1, 1'b1, 0, 0) c177052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177052));
	wire w193052;
	repeater #(1, 1'b1, 0, 0) c193052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193052));
	wire w3053;
	repeater #(1, 1'b1, 0, 0) c3053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3053));
	wire w19053;
	repeater #(1, 1'b1, 0, 0) c19053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19053));
	wire w73053;
	assign outputs[15] = ();
	wire w133053;
	repeater #(1, 1'b0, 0, 0) c133053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133053));
	wire w190054;
	torch #(1'b1) c190054 (.i_clk(tick), .i_in(), .o_out(w190054));
	wire w16055;
	torch #(1'b1) c16055 (.i_clk(tick), .i_in(), .o_out(w16055));
	wire w103055;
	repeater #(1, 1'b0, 0, 0) c103055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103055));
	wire w182056;
	torch #(1'b1) c182056 (.i_clk(tick), .i_in(), .o_out(w182056));
	wire w198056;
	torch #(1'b1) c198056 (.i_clk(tick), .i_in(), .o_out(w198056));
	wire w8057;
	torch #(1'b1) c8057 (.i_clk(tick), .i_in(), .o_out(w8057));
	wire w24057;
	torch #(1'b1) c24057 (.i_clk(tick), .i_in(), .o_out(w24057));
	wire w189057;
	repeater #(1, 1'b0, 0, 0) c189057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189057));
	wire w15058;
	repeater #(1, 1'b0, 0, 0) c15058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15058));
	wire w112058;
	torch #(1'b1) c112058 (.i_clk(tick), .i_in(), .o_out(w112058));
	wire w116058;
	torch #(1'b1) c116058 (.i_clk(tick), .i_in(), .o_out(w116058));
	wire w120058;
	torch #(1'b1) c120058 (.i_clk(tick), .i_in(), .o_out(w120058));
	wire w124058;
	torch #(1'b1) c124058 (.i_clk(tick), .i_in(), .o_out(w124058));
	wire w183058;
	repeater #(1, 1'b0, 0, 0) c183058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183058));
	wire w199058;
	repeater #(1, 1'b0, 0, 0) c199058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199058));
	wire w9059;
	repeater #(1, 1'b0, 0, 0) c9059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9059));
	wire w25059;
	repeater #(1, 1'b0, 0, 0) c25059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25059));
	wire w105062;
	torch #(1'b0) c105062 (.i_clk(tick), .i_in(), .o_out(w105062));
	wire w109062;
	torch #(1'b0) c109062 (.i_clk(tick), .i_in(), .o_out(w109062));
	wire w113062;
	torch #(1'b0) c113062 (.i_clk(tick), .i_in(), .o_out(w113062));
	wire w117062;
	torch #(1'b0) c117062 (.i_clk(tick), .i_in(), .o_out(w117062));
	wire w121062;
	torch #(1'b0) c121062 (.i_clk(tick), .i_in(), .o_out(w121062));
	wire w125062;
	torch #(1'b0) c125062 (.i_clk(tick), .i_in(), .o_out(w125062));
	wire w129062;
	torch #(1'b0) c129062 (.i_clk(tick), .i_in(), .o_out(w129062));
	wire w106064;
	torch #(1'b1) c106064 (.i_clk(tick), .i_in(), .o_out(w106064));
	wire w110064;
	torch #(1'b1) c110064 (.i_clk(tick), .i_in(), .o_out(w110064));
	wire w114064;
	torch #(1'b1) c114064 (.i_clk(tick), .i_in(), .o_out(w114064));
	wire w118064;
	torch #(1'b1) c118064 (.i_clk(tick), .i_in(), .o_out(w118064));
	wire w122064;
	torch #(1'b1) c122064 (.i_clk(tick), .i_in(), .o_out(w122064));
	wire w126064;
	torch #(1'b1) c126064 (.i_clk(tick), .i_in(), .o_out(w126064));
	wire w130064;
	torch #(1'b1) c130064 (.i_clk(tick), .i_in(), .o_out(w130064));
	wire w107066;
	torch #(1'b0) c107066 (.i_clk(tick), .i_in(), .o_out(w107066));
	wire w111066;
	torch #(1'b0) c111066 (.i_clk(tick), .i_in(), .o_out(w111066));
	wire w115066;
	torch #(1'b0) c115066 (.i_clk(tick), .i_in(), .o_out(w115066));
	wire w119066;
	torch #(1'b0) c119066 (.i_clk(tick), .i_in(), .o_out(w119066));
	wire w123066;
	torch #(1'b0) c123066 (.i_clk(tick), .i_in(), .o_out(w123066));
	wire w127066;
	torch #(1'b0) c127066 (.i_clk(tick), .i_in(), .o_out(w127066));
	wire w131066;
	torch #(1'b0) c131066 (.i_clk(tick), .i_in(), .o_out(w131066));
	wire w133069;
	repeater #(1, 1'b0, 0, 0) c133069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133069));
	wire w103071;
	repeater #(1, 1'b0, 0, 0) c103071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103071));
	wire w112074;
	torch #(1'b1) c112074 (.i_clk(tick), .i_in(), .o_out(w112074));
	wire w116074;
	torch #(1'b1) c116074 (.i_clk(tick), .i_in(), .o_out(w116074));
	wire w120074;
	torch #(1'b1) c120074 (.i_clk(tick), .i_in(), .o_out(w120074));
	wire w124074;
	torch #(1'b1) c124074 (.i_clk(tick), .i_in(), .o_out(w124074));
	wire w60075;

	wire w78075;

	wire w105078;
	torch #(1'b0) c105078 (.i_clk(tick), .i_in(), .o_out(w105078));
	wire w109078;
	torch #(1'b0) c109078 (.i_clk(tick), .i_in(), .o_out(w109078));
	wire w113078;
	torch #(1'b0) c113078 (.i_clk(tick), .i_in(), .o_out(w113078));
	wire w117078;
	torch #(1'b1) c117078 (.i_clk(tick), .i_in(), .o_out(w117078));
	wire w121078;
	torch #(1'b0) c121078 (.i_clk(tick), .i_in(), .o_out(w121078));
	wire w125078;
	torch #(1'b0) c125078 (.i_clk(tick), .i_in(), .o_out(w125078));
	wire w129078;
	torch #(1'b0) c129078 (.i_clk(tick), .i_in(), .o_out(w129078));
	wire w106080;
	torch #(1'b1) c106080 (.i_clk(tick), .i_in(), .o_out(w106080));
	wire w110080;
	torch #(1'b1) c110080 (.i_clk(tick), .i_in(), .o_out(w110080));
	wire w114080;
	torch #(1'b1) c114080 (.i_clk(tick), .i_in(), .o_out(w114080));
	wire w118080;
	torch #(1'b1) c118080 (.i_clk(tick), .i_in(), .o_out(w118080));
	wire w122080;
	torch #(1'b1) c122080 (.i_clk(tick), .i_in(), .o_out(w122080));
	wire w126080;
	torch #(1'b1) c126080 (.i_clk(tick), .i_in(), .o_out(w126080));
	wire w130080;
	torch #(1'b1) c130080 (.i_clk(tick), .i_in(), .o_out(w130080));
	wire w107082;
	torch #(1'b0) c107082 (.i_clk(tick), .i_in(), .o_out(w107082));
	wire w111082;
	torch #(1'b0) c111082 (.i_clk(tick), .i_in(), .o_out(w111082));
	wire w115082;
	torch #(1'b0) c115082 (.i_clk(tick), .i_in(), .o_out(w115082));
	wire w119082;
	torch #(1'b0) c119082 (.i_clk(tick), .i_in(), .o_out(w119082));
	wire w123082;
	torch #(1'b0) c123082 (.i_clk(tick), .i_in(), .o_out(w123082));
	wire w127082;
	torch #(1'b0) c127082 (.i_clk(tick), .i_in(), .o_out(w127082));
	wire w131082;
	torch #(1'b0) c131082 (.i_clk(tick), .i_in(), .o_out(w131082));
	wire w133085;
	repeater #(1, 1'b0, 0, 0) c133085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133085));
	wire w103087;
	repeater #(1, 1'b0, 0, 0) c103087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103087));
	wire w112090;
	torch #(1'b1) c112090 (.i_clk(tick), .i_in(), .o_out(w112090));
	wire w116090;
	torch #(1'b1) c116090 (.i_clk(tick), .i_in(), .o_out(w116090));
	wire w120090;
	torch #(1'b1) c120090 (.i_clk(tick), .i_in(), .o_out(w120090));
	wire w124090;
	torch #(1'b1) c124090 (.i_clk(tick), .i_in(), .o_out(w124090));
	wire w105094;
	torch #(1'b0) c105094 (.i_clk(tick), .i_in(), .o_out(w105094));
	wire w109094;
	torch #(1'b0) c109094 (.i_clk(tick), .i_in(), .o_out(w109094));
	wire w113094;
	torch #(1'b0) c113094 (.i_clk(tick), .i_in(), .o_out(w113094));
	wire w117094;
	torch #(1'b0) c117094 (.i_clk(tick), .i_in(), .o_out(w117094));
	wire w121094;
	torch #(1'b0) c121094 (.i_clk(tick), .i_in(), .o_out(w121094));
	wire w125094;
	torch #(1'b0) c125094 (.i_clk(tick), .i_in(), .o_out(w125094));
	wire w129094;
	torch #(1'b0) c129094 (.i_clk(tick), .i_in(), .o_out(w129094));
	wire w106096;
	torch #(1'b1) c106096 (.i_clk(tick), .i_in(), .o_out(w106096));
	wire w110096;
	torch #(1'b1) c110096 (.i_clk(tick), .i_in(), .o_out(w110096));
	wire w114096;
	torch #(1'b1) c114096 (.i_clk(tick), .i_in(), .o_out(w114096));
	wire w118096;
	torch #(1'b1) c118096 (.i_clk(tick), .i_in(), .o_out(w118096));
	wire w122096;
	torch #(1'b1) c122096 (.i_clk(tick), .i_in(), .o_out(w122096));
	wire w126096;
	torch #(1'b1) c126096 (.i_clk(tick), .i_in(), .o_out(w126096));
	wire w130096;
	torch #(1'b1) c130096 (.i_clk(tick), .i_in(), .o_out(w130096));
	wire w107098;
	torch #(1'b0) c107098 (.i_clk(tick), .i_in(), .o_out(w107098));
	wire w111098;
	torch #(1'b0) c111098 (.i_clk(tick), .i_in(), .o_out(w111098));
	wire w115098;
	torch #(1'b0) c115098 (.i_clk(tick), .i_in(), .o_out(w115098));
	wire w119098;
	torch #(1'b0) c119098 (.i_clk(tick), .i_in(), .o_out(w119098));
	wire w123098;
	torch #(1'b0) c123098 (.i_clk(tick), .i_in(), .o_out(w123098));
	wire w127098;
	torch #(1'b0) c127098 (.i_clk(tick), .i_in(), .o_out(w127098));
	wire w131098;
	torch #(1'b0) c131098 (.i_clk(tick), .i_in(), .o_out(w131098));
	wire w1030108;
	repeater #(2, 1'b0, 0, 0) c1030108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030108));
	wire w1070108;
	repeater #(2, 1'b0, 0, 0) c1070108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070108));
	wire w1110108;
	repeater #(2, 1'b0, 0, 0) c1110108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110108));
	wire w1150108;
	repeater #(2, 1'b0, 0, 0) c1150108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1150108));
	wire w1190108;
	repeater #(2, 1'b0, 0, 0) c1190108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190108));
	wire w1230108;
	repeater #(2, 1'b0, 0, 0) c1230108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230108));
	wire w1270108;
	repeater #(2, 1'b0, 0, 0) c1270108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1270108));
	wire w1040110;

	wire w1080110;

	wire w1120110;

	wire w1160110;

	wire w1200110;

	wire w1240110;

	wire w1280110;

	wire w1040111;

	wire w1080111;

	wire w1120111;

	wire w1160111;

	wire w1200111;

	wire w1240111;

	wire w1280111;

	wire w1030114;
	repeater #(1, 1'b1, 0, 0) c1030114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030114));
	wire w1070114;
	repeater #(1, 1'b1, 0, 0) c1070114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070114));
	wire w1110114;
	repeater #(1, 1'b1, 0, 0) c1110114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110114));
	wire w1150114;
	repeater #(1, 1'b0, 0, 0) c1150114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1150114));
	wire w1190114;
	repeater #(1, 1'b1, 0, 0) c1190114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190114));
	wire w1230114;
	repeater #(1, 1'b1, 0, 0) c1230114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230114));
	wire w1270114;
	repeater #(1, 1'b1, 0, 0) c1270114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1270114));
	wire w1050115;

	wire w1090115;

	wire w1130115;

	wire w1170115;

	wire w1210115;

	wire w1250115;

	wire w1290115;

	wire w1040116;

	wire w1080116;

	wire w1120116;

	wire w1160116;

	wire w1200116;

	wire w1240116;

	wire w1280116;

	wire w1060118;
	torch #(1'b0) c1060118 (.i_clk(tick), .i_in(), .o_out(w1060118));
	wire w1100118;
	torch #(1'b0) c1100118 (.i_clk(tick), .i_in(), .o_out(w1100118));
	wire w1140118;
	torch #(1'b1) c1140118 (.i_clk(tick), .i_in(), .o_out(w1140118));
	wire w1180118;
	torch #(1'b1) c1180118 (.i_clk(tick), .i_in(), .o_out(w1180118));
	wire w1220118;
	torch #(1'b1) c1220118 (.i_clk(tick), .i_in(), .o_out(w1220118));
	wire w1260118;
	torch #(1'b0) c1260118 (.i_clk(tick), .i_in(), .o_out(w1260118));
	wire w1300118;
	torch #(1'b0) c1300118 (.i_clk(tick), .i_in(), .o_out(w1300118));
	wire w1030119;
	torch #(1'b0) c1030119 (.i_clk(tick), .i_in(), .o_out(w1030119));
	wire w1050119;
	torch #(1'b0) c1050119 (.i_clk(tick), .i_in(), .o_out(w1050119));
	wire w1070119;
	torch #(1'b0) c1070119 (.i_clk(tick), .i_in(), .o_out(w1070119));
	wire w1090119;
	torch #(1'b0) c1090119 (.i_clk(tick), .i_in(), .o_out(w1090119));
	wire w1110119;
	torch #(1'b0) c1110119 (.i_clk(tick), .i_in(), .o_out(w1110119));
	wire w1130119;
	torch #(1'b0) c1130119 (.i_clk(tick), .i_in(), .o_out(w1130119));
	wire w1150119;
	torch #(1'b0) c1150119 (.i_clk(tick), .i_in(), .o_out(w1150119));
	wire w1170119;
	torch #(1'b0) c1170119 (.i_clk(tick), .i_in(), .o_out(w1170119));
	wire w1190119;
	torch #(1'b0) c1190119 (.i_clk(tick), .i_in(), .o_out(w1190119));
	wire w1210119;
	torch #(1'b0) c1210119 (.i_clk(tick), .i_in(), .o_out(w1210119));
	wire w1230119;
	torch #(1'b0) c1230119 (.i_clk(tick), .i_in(), .o_out(w1230119));
	wire w1250119;
	torch #(1'b0) c1250119 (.i_clk(tick), .i_in(), .o_out(w1250119));
	wire w1270119;
	torch #(1'b0) c1270119 (.i_clk(tick), .i_in(), .o_out(w1270119));
	wire w1290119;
	torch #(1'b0) c1290119 (.i_clk(tick), .i_in(), .o_out(w1290119));
	wire w2020156;

	wire w270157;

	wire w280157;

	wire w610157;

	wire w620157;

	wire w950157;

	wire w960157;

	wire w1290157;

	wire w2030157;
	repeater #(1, 1'b1, 0, 0) c2030157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030157));
	wire w290158;
	repeater #(1, 1'b1, 0, 0) c290158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290158));
	wire w630158;
	repeater #(1, 1'b1, 0, 0) c630158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630158));
	wire w970158;
	repeater #(1, 1'b1, 0, 0) c970158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w970158));
	wire w2000158;

	wire w250159;

	wire w260159;

	wire w590159;

	wire w600159;

	wire w930159;

	wire w940159;

	wire w1270159;

	wire w1300159;
	repeater #(1, 1'b1, 0, 0) c1300159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1300159));
	wire w2010159;
	repeater #(1, 1'b1, 0, 0) c2010159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010159));
	wire w270160;
	repeater #(1, 1'b1, 0, 0) c270160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w270160));
	wire w610160;
	repeater #(1, 1'b1, 0, 0) c610160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w610160));
	wire w950160;
	repeater #(1, 1'b1, 0, 0) c950160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w950160));
	wire w1290160;

	wire w1980160;

	wire w230161;

	wire w240161;

	wire w570161;

	wire w580161;

	wire w910161;

	wire w920161;

	wire w1250161;

	wire w1280161;
	repeater #(1, 1'b1, 0, 0) c1280161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1280161));
	wire w1990161;
	repeater #(1, 1'b1, 0, 0) c1990161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990161));
	wire w250162;
	repeater #(1, 1'b1, 0, 0) c250162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250162));
	wire w590162;
	repeater #(1, 1'b1, 0, 0) c590162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590162));
	wire w930162;
	repeater #(1, 1'b1, 0, 0) c930162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w930162));
	wire w1270162;

	wire w1960162;

	wire w210163;

	wire w220163;

	wire w550163;

	wire w560163;

	wire w890163;

	wire w900163;

	wire w1230163;

	wire w1260163;
	repeater #(1, 1'b1, 0, 0) c1260163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1260163));
	wire w1970163;
	repeater #(1, 1'b1, 0, 0) c1970163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970163));
	wire w230164;
	repeater #(1, 1'b1, 0, 0) c230164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230164));
	wire w570164;
	repeater #(1, 1'b1, 0, 0) c570164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570164));
	wire w910164;
	repeater #(1, 1'b1, 0, 0) c910164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w910164));
	wire w1250164;

	wire w1940164;

	wire w190165;

	wire w200165;

	wire w530165;

	wire w540165;

	wire w870165;

	wire w880165;

	wire w1210165;

	wire w1240165;
	repeater #(1, 1'b1, 0, 0) c1240165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240165));
	wire w1950165;
	repeater #(1, 1'b1, 0, 0) c1950165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950165));
	wire w210166;
	repeater #(1, 1'b1, 0, 0) c210166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210166));
	wire w550166;
	repeater #(1, 1'b1, 0, 0) c550166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550166));
	wire w890166;
	repeater #(1, 1'b1, 0, 0) c890166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w890166));
	wire w1230166;

	wire w1920166;

	wire w170167;

	wire w180167;

	wire w510167;

	wire w520167;

	wire w850167;

	wire w860167;

	wire w1190167;

	wire w1220167;
	repeater #(1, 1'b1, 0, 0) c1220167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1220167));
	wire w1930167;
	repeater #(1, 1'b1, 0, 0) c1930167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1930167));
	wire w190168;
	repeater #(1, 1'b1, 0, 0) c190168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190168));
	wire w530168;
	repeater #(1, 1'b1, 0, 0) c530168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530168));
	wire w870168;
	repeater #(1, 1'b1, 0, 0) c870168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w870168));
	wire w1210168;

	wire w1900168;

	wire w150169;

	wire w160169;

	wire w490169;

	wire w500169;

	wire w830169;

	wire w840169;

	wire w1170169;

	wire w1200169;
	repeater #(1, 1'b1, 0, 0) c1200169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1200169));
	wire w1910169;
	repeater #(1, 1'b0, 0, 0) c1910169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910169));
	wire w170170;
	repeater #(1, 1'b0, 0, 0) c170170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170170));
	wire w510170;
	repeater #(1, 1'b0, 0, 0) c510170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510170));
	wire w850170;
	repeater #(1, 1'b0, 0, 0) c850170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w850170));
	wire w1190170;

	wire w1880170;

	wire w130171;

	wire w140171;

	wire w470171;

	wire w480171;

	wire w810171;

	wire w820171;

	wire w1150171;

	wire w1180171;
	repeater #(1, 1'b0, 0, 0) c1180171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1180171));
	wire w1890171;
	repeater #(1, 1'b0, 0, 0) c1890171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1890171));
	wire w150172;
	repeater #(1, 1'b0, 0, 0) c150172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150172));
	wire w490172;
	repeater #(1, 1'b0, 0, 0) c490172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w490172));
	wire w830172;
	repeater #(1, 1'b0, 0, 0) c830172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w830172));
	wire w1170172;

	wire w1860172;

	wire w110173;

	wire w120173;

	wire w450173;

	wire w460173;

	wire w790173;

	wire w800173;

	wire w1130173;

	wire w1160173;
	repeater #(1, 1'b0, 0, 0) c1160173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1160173));
	wire w1870173;
	repeater #(1, 1'b1, 0, 0) c1870173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870173));
	wire w130174;
	repeater #(1, 1'b1, 0, 0) c130174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130174));
	wire w470174;
	repeater #(1, 1'b1, 0, 0) c470174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470174));
	wire w810174;
	repeater #(1, 1'b1, 0, 0) c810174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w810174));
	wire w1150174;

	wire w1840174;

	wire w90175;

	wire w100175;

	wire w430175;

	wire w440175;

	wire w770175;

	wire w780175;

	wire w1110175;

	wire w1140175;
	repeater #(1, 1'b1, 0, 0) c1140175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1140175));
	wire w1850175;
	repeater #(1, 1'b1, 0, 0) c1850175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850175));
	wire w110176;
	repeater #(1, 1'b1, 0, 0) c110176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110176));
	wire w450176;
	repeater #(1, 1'b1, 0, 0) c450176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w450176));
	wire w790176;
	repeater #(1, 1'b1, 0, 0) c790176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w790176));
	wire w1130176;

	wire w1820176;

	wire w70177;

	wire w80177;

	wire w410177;

	wire w420177;

	wire w750177;

	wire w760177;

	wire w1090177;

	wire w1120177;
	repeater #(1, 1'b1, 0, 0) c1120177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1120177));
	wire w1830177;
	repeater #(1, 1'b1, 0, 0) c1830177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830177));
	wire w90178;
	repeater #(1, 1'b1, 0, 0) c90178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90178));
	wire w430178;
	repeater #(1, 1'b1, 0, 0) c430178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w430178));
	wire w770178;
	repeater #(1, 1'b1, 0, 0) c770178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w770178));
	wire w1110178;

	wire w1800178;

	wire w510;

	wire w610;

	wire w3910;

	wire w4010;

	wire w7310;

	wire w7410;

	wire w10710;

	wire w11010;
	repeater #(1, 1'b1, 0, 0) c11010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11010));
	wire w18110;
	repeater #(1, 1'b1, 0, 0) c18110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18110));
	wire w711;
	repeater #(1, 1'b1, 0, 0) c711 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711));
	wire w4111;
	repeater #(1, 1'b1, 0, 0) c4111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4111));
	wire w7511;
	repeater #(1, 1'b1, 0, 0) c7511 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7511));
	wire w10911;

	wire w17811;

	wire w312;

	wire w412;

	wire w3712;

	wire w3812;

	wire w7112;

	wire w7212;

	wire w10512;

	wire w10812;
	repeater #(1, 1'b1, 0, 0) c10812 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10812));
	wire w17912;
	repeater #(1, 1'b1, 0, 0) c17912 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17912));
	wire w513;
	repeater #(1, 1'b1, 0, 0) c513 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w513));
	wire w3913;
	repeater #(1, 1'b1, 0, 0) c3913 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3913));
	wire w7313;
	repeater #(1, 1'b1, 0, 0) c7313 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7313));
	wire w10713;

	wire w114;

	wire w3514;

	wire w6914;

	wire w10314;

	wire w10614;
	repeater #(1, 1'b1, 0, 0) c10614 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10614));
	wire w17714;
	repeater #(1, 1'b1, 0, 0) c17714 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17714));
	wire w315;
	repeater #(1, 1'b1, 0, 0) c315 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w315));
	wire w3715;
	repeater #(1, 1'b1, 0, 0) c3715 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3715));
	wire w7115;
	repeater #(1, 1'b1, 0, 0) c7115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7115));
	wire w10515;

	wire w10416;
	repeater #(2, 1'b1, 0, 0) c10416 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10416));
	wire w10617;
	repeater #(1, 1'b1, 0, 0) c10617 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10617));
	wire w19619;
	repeater #(2, 1'b1, 0, 0) c19619 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19619));
	wire w22110;
	repeater #(2, 1'b1, 0, 0) c22110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22110));
	wire w105110;
	torch #(1'b1) c105110 (.i_clk(tick), .i_in(), .o_out(w105110));
	wire w109110;
	torch #(1'b1) c109110 (.i_clk(tick), .i_in(), .o_out(w109110));
	wire w113110;
	torch #(1'b1) c113110 (.i_clk(tick), .i_in(), .o_out(w113110));
	wire w117110;
	torch #(1'b1) c117110 (.i_clk(tick), .i_in(), .o_out(w117110));
	wire w121110;
	torch #(1'b1) c121110 (.i_clk(tick), .i_in(), .o_out(w121110));
	wire w125110;
	torch #(1'b1) c125110 (.i_clk(tick), .i_in(), .o_out(w125110));
	wire w129110;
	torch #(1'b1) c129110 (.i_clk(tick), .i_in(), .o_out(w129110));
	wire w182111;
	repeater #(1, 1'b1, 0, 0) c182111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182111));
	wire w188111;
	torch #(1'b0) c188111 (.i_clk(tick), .i_in(), .o_out(w188111));
	wire w198111;
	repeater #(1, 1'b1, 0, 0) c198111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198111));
	wire w8112;
	repeater #(1, 1'b1, 0, 0) c8112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8112));
	wire w14112;
	torch #(1'b0) c14112 (.i_clk(tick), .i_in(), .o_out(w14112));
	wire w24112;
	repeater #(1, 1'b1, 0, 0) c24112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24112));
	wire w106113;
	repeater #(1, 1'b1, 0, 0) c106113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106113));
	wire w110113;
	repeater #(1, 1'b1, 0, 0) c110113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110113));
	wire w114113;
	repeater #(1, 1'b1, 0, 0) c114113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114113));
	wire w118113;
	repeater #(1, 1'b1, 0, 0) c118113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118113));
	wire w122113;
	repeater #(1, 1'b1, 0, 0) c122113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122113));
	wire w126113;
	repeater #(1, 1'b1, 0, 0) c126113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126113));
	wire w130113;
	repeater #(1, 1'b1, 0, 0) c130113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130113));
	wire w105114;
	torch #(1'b1) c105114 (.i_clk(tick), .i_in(), .o_out(w105114));
	wire w109114;
	torch #(1'b1) c109114 (.i_clk(tick), .i_in(), .o_out(w109114));
	wire w113114;
	torch #(1'b1) c113114 (.i_clk(tick), .i_in(), .o_out(w113114));
	wire w117114;
	torch #(1'b1) c117114 (.i_clk(tick), .i_in(), .o_out(w117114));
	wire w121114;
	torch #(1'b1) c121114 (.i_clk(tick), .i_in(), .o_out(w121114));
	wire w125114;
	torch #(1'b1) c125114 (.i_clk(tick), .i_in(), .o_out(w125114));
	wire w129114;
	torch #(1'b1) c129114 (.i_clk(tick), .i_in(), .o_out(w129114));
	wire w189114;
	repeater #(1, 1'b0, 0, 0) c189114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189114));
	wire w15115;
	repeater #(1, 1'b1, 0, 0) c15115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15115));
	wire w182115;
	repeater #(1, 1'b1, 0, 0) c182115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182115));
	wire w198115;
	repeater #(1, 1'b1, 0, 0) c198115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198115));
	wire w8116;
	repeater #(1, 1'b1, 0, 0) c8116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8116));
	wire w24116;
	repeater #(1, 1'b1, 0, 0) c24116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24116));
	wire w43116;
	torch #(1'b1) c43116 (.i_clk(tick), .i_in(), .o_out(w43116));
	wire w47116;
	torch #(1'b0) c47116 (.i_clk(tick), .i_in(), .o_out(w47116));
	wire w51116;
	torch #(1'b1) c51116 (.i_clk(tick), .i_in(), .o_out(w51116));
	wire w55116;
	torch #(1'b1) c55116 (.i_clk(tick), .i_in(), .o_out(w55116));
	wire w79116;
	torch #(1'b0) c79116 (.i_clk(tick), .i_in(), .o_out(w79116));
	wire w83116;
	torch #(1'b0) c83116 (.i_clk(tick), .i_in(), .o_out(w83116));
	wire w87116;
	torch #(1'b1) c87116 (.i_clk(tick), .i_in(), .o_out(w87116));
	wire w91116;
	torch #(1'b0) c91116 (.i_clk(tick), .i_in(), .o_out(w91116));
	wire w187116;

	wire w13117;

	wire w104117;
	torch #(1'b0) c104117 (.i_clk(tick), .i_in(), .o_out(w104117));
	wire w108117;
	torch #(1'b0) c108117 (.i_clk(tick), .i_in(), .o_out(w108117));
	wire w112117;
	torch #(1'b0) c112117 (.i_clk(tick), .i_in(), .o_out(w112117));
	wire w116117;
	torch #(1'b1) c116117 (.i_clk(tick), .i_in(), .o_out(w116117));
	wire w120117;
	torch #(1'b0) c120117 (.i_clk(tick), .i_in(), .o_out(w120117));
	wire w124117;
	torch #(1'b0) c124117 (.i_clk(tick), .i_in(), .o_out(w124117));
	wire w128117;
	torch #(1'b0) c128117 (.i_clk(tick), .i_in(), .o_out(w128117));
	wire w179117;

	wire w195117;

	wire w5118;

	wire w21118;

	wire w176118;

	wire w181118;

	wire w182118;

	wire w192118;

	wire w197118;

	wire w198118;

	wire w2119;

	wire w7119;

	wire w8119;

	wire w18119;

	wire w23119;

	wire w24119;

	wire w174120;

	wire w190120;

	wire w0121;

	wire w16121;

	wire w180121;

	wire w181121;

	wire w196121;

	wire w197121;

	wire w6122;

	wire w7122;

	wire w22122;

	wire w23122;

	wire w190122;

	wire w16123;

	wire w43123;
	repeater #(2, 1'b0, 0, 0) c43123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43123));
	wire w45123;
	repeater #(1, 1'b0, 0, 0) c45123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45123));
	wire w47123;
	repeater #(2, 1'b1, 0, 0) c47123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47123));
	wire w49123;
	repeater #(1, 1'b0, 0, 0) c49123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49123));
	wire w51123;
	repeater #(2, 1'b0, 0, 0) c51123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51123));
	wire w53123;
	repeater #(1, 1'b0, 0, 0) c53123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53123));
	wire w55123;
	repeater #(2, 1'b0, 0, 0) c55123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55123));
	wire w57123;
	repeater #(1, 1'b0, 0, 0) c57123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57123));
	wire w77123;
	repeater #(1, 1'b1, 0, 0) c77123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77123));
	wire w79123;
	repeater #(2, 1'b1, 0, 0) c79123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79123));
	wire w81123;
	repeater #(1, 1'b1, 0, 0) c81123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81123));
	wire w83123;
	repeater #(2, 1'b1, 0, 0) c83123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83123));
	wire w85123;
	repeater #(1, 1'b1, 0, 0) c85123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85123));
	wire w87123;
	repeater #(2, 1'b0, 0, 0) c87123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87123));
	wire w89123;
	repeater #(1, 1'b1, 0, 0) c89123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89123));
	wire w91123;
	repeater #(2, 1'b1, 0, 0) c91123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91123));
	wire w112123;
	torch #(1'b1) c112123 (.i_clk(tick), .i_in(), .o_out(w112123));
	wire w116123;
	torch #(1'b1) c116123 (.i_clk(tick), .i_in(), .o_out(w116123));
	wire w120123;
	torch #(1'b1) c120123 (.i_clk(tick), .i_in(), .o_out(w120123));
	wire w124123;
	torch #(1'b1) c124123 (.i_clk(tick), .i_in(), .o_out(w124123));
	wire w174124;

	wire w178124;

	wire w182124;

	wire w186124;

	wire w190124;

	wire w194124;

	wire w198124;

	wire w0125;

	wire w4125;

	wire w8125;

	wire w12125;

	wire w16125;

	wire w20125;

	wire w24125;

	wire w52125;

	wire w82125;

	wire w44126;

	wire w48126;

	wire w51126;

	wire w53126;

	wire w56126;

	wire w78126;

	wire w81126;

	wire w83126;

	wire w86126;

	wire w90126;

	wire w43127;

	wire w45127;

	wire w47127;

	wire w49127;

	wire w52127;

	wire w55127;

	wire w57127;

	wire w77127;

	wire w79127;

	wire w82127;

	wire w85127;

	wire w87127;

	wire w89127;

	wire w91127;

	wire w48128;

	wire w86128;

	wire w174128;

	wire w178128;

	wire w182128;

	wire w186128;

	wire w190128;

	wire w194128;

	wire w198128;

	wire w0129;

	wire w4129;

	wire w8129;

	wire w12129;

	wire w16129;

	wire w20129;

	wire w24129;

	wire w44129;

	wire w48129;

	wire w49129;

	wire w53129;

	wire w55129;

	wire w57129;

	wire w77129;

	wire w79129;

	wire w81129;

	wire w85129;

	wire w86129;

	wire w90129;

	wire w48130;

	wire w86130;

	wire w172130;
	repeater #(1, 1'b1, 0, 0) c172130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172130));
	wire w176130;
	repeater #(1, 1'b1, 0, 0) c176130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176130));
	wire w180130;
	repeater #(1, 1'b1, 0, 0) c180130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180130));
	wire w184130;
	repeater #(1, 1'b0, 0, 0) c184130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184130));
	wire w206130;
	repeater #(1, 1'b1, 0, 0) c206130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206130));
	wire w2131;
	repeater #(1, 1'b1, 0, 0) c2131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2131));
	wire w6131;
	repeater #(1, 1'b1, 0, 0) c6131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6131));
	wire w10131;
	repeater #(1, 1'b1, 0, 0) c10131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10131));
	wire w41131;

	wire w46131;

	wire w47131;

	wire w87131;

	wire w88131;

	wire w93131;

	wire w190131;

	wire w194131;

	wire w198131;

	wire w16132;

	wire w20132;

	wire w24132;

	wire w39132;
	repeater #(1, 1'b1, 0, 0) c39132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39132));
	wire w44132;
	repeater #(1, 1'b1, 0, 0) c44132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44132));
	wire w90132;
	repeater #(1, 1'b1, 0, 0) c90132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90132));
	wire w95132;
	repeater #(1, 1'b1, 0, 0) c95132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95132));
	wire w105132;
	torch #(1'b1) c105132 (.i_clk(tick), .i_in(), .o_out(w105132));
	wire w109132;
	torch #(1'b1) c109132 (.i_clk(tick), .i_in(), .o_out(w109132));
	wire w113132;
	torch #(1'b1) c113132 (.i_clk(tick), .i_in(), .o_out(w113132));
	wire w117132;
	torch #(1'b1) c117132 (.i_clk(tick), .i_in(), .o_out(w117132));
	wire w121132;
	torch #(1'b1) c121132 (.i_clk(tick), .i_in(), .o_out(w121132));
	wire w125132;
	torch #(1'b1) c125132 (.i_clk(tick), .i_in(), .o_out(w125132));
	wire w129132;
	torch #(1'b1) c129132 (.i_clk(tick), .i_in(), .o_out(w129132));
	wire w49133;
	repeater #(1, 1'b1, 0, 0) c49133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49133));
	wire w85133;
	repeater #(1, 1'b0, 0, 0) c85133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85133));
	wire w106133;
	repeater #(1, 1'b0, 0, 0) c106133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106133));
	wire w110133;
	repeater #(1, 1'b0, 0, 0) c110133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110133));
	wire w114133;
	repeater #(1, 1'b0, 0, 0) c114133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114133));
	wire w118133;
	repeater #(1, 1'b1, 0, 0) c118133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118133));
	wire w122133;
	repeater #(1, 1'b0, 0, 0) c122133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122133));
	wire w126133;
	repeater #(1, 1'b0, 0, 0) c126133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126133));
	wire w130133;
	repeater #(1, 1'b0, 0, 0) c130133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130133));
	wire w190133;

	wire w16134;

	wire w172134;
	repeater #(1, 1'b1, 0, 0) c172134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172134));
	wire w188134;
	repeater #(1, 1'b1, 0, 0) c188134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188134));
	wire w206134;
	repeater #(1, 1'b1, 0, 0) c206134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206134));
	wire w14135;
	repeater #(1, 1'b1, 0, 0) c14135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14135));
	wire w104135;

	wire w106135;
	repeater #(1, 1'b0, 0, 0) c106135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106135));
	wire w108135;

	wire w110135;
	repeater #(1, 1'b0, 0, 0) c110135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110135));
	wire w112135;

	wire w114135;
	repeater #(1, 1'b0, 0, 0) c114135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114135));
	wire w116135;

	wire w118135;
	repeater #(1, 1'b1, 0, 0) c118135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118135));
	wire w120135;

	wire w122135;
	repeater #(1, 1'b0, 0, 0) c122135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122135));
	wire w124135;

	wire w126135;
	repeater #(1, 1'b0, 0, 0) c126135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126135));
	wire w128135;

	wire w130135;
	repeater #(1, 1'b0, 0, 0) c130135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130135));
	wire w179135;
	repeater #(1, 1'b1, 0, 0) c179135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179135));
	wire w195135;
	repeater #(1, 1'b1, 0, 0) c195135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195135));
	wire w5136;
	repeater #(1, 1'b1, 0, 0) c5136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5136));
	wire w21136;
	repeater #(1, 1'b1, 0, 0) c21136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21136));
	wire w39136;
	repeater #(1, 1'b1, 0, 0) c39136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39136));
	wire w44136;
	repeater #(1, 1'b0, 0, 0) c44136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44136));
	wire w49136;
	repeater #(1, 1'b0, 0, 0) c49136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49136));
	wire w85136;
	repeater #(1, 1'b0, 0, 0) c85136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85136));
	wire w90136;
	repeater #(1, 1'b1, 0, 0) c90136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90136));
	wire w95136;
	repeater #(1, 1'b1, 0, 0) c95136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95136));
	wire w174136;

	wire w190136;

	wire w0137;

	wire w16137;

	wire w182137;

	wire w8138;

	wire w177138;

	wire w179138;

	wire w180138;

	wire w185138;

	wire w193138;

	wire w195138;

	wire w196138;

	wire w3139;

	wire w5139;

	wire w6139;

	wire w11139;

	wire w19139;

	wire w21139;

	wire w22139;

	wire w112139;
	torch #(1'b1) c112139 (.i_clk(tick), .i_in(), .o_out(w112139));
	wire w116139;
	torch #(1'b1) c116139 (.i_clk(tick), .i_in(), .o_out(w116139));
	wire w120139;
	torch #(1'b1) c120139 (.i_clk(tick), .i_in(), .o_out(w120139));
	wire w124139;
	torch #(1'b1) c124139 (.i_clk(tick), .i_in(), .o_out(w124139));
	wire w39140;
	repeater #(1, 1'b0, 0, 0) c39140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39140));
	wire w44140;
	repeater #(1, 1'b0, 0, 0) c44140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44140));
	wire w49140;
	repeater #(1, 1'b0, 0, 0) c49140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49140));
	wire w85140;
	repeater #(1, 1'b0, 0, 0) c85140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85140));
	wire w90140;
	repeater #(1, 1'b1, 0, 0) c90140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90140));
	wire w95140;
	repeater #(1, 1'b1, 0, 0) c95140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95140));
	wire w187140;

	wire w188140;

	wire w13141;

	wire w14141;

	wire w177142;

	wire w179142;

	wire w180142;

	wire w193142;

	wire w195142;

	wire w196142;

	wire w3143;

	wire w5143;

	wire w6143;

	wire w19143;

	wire w21143;

	wire w22143;

	wire w39144;
	repeater #(2, 1'b0, 0, 0) c39144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39144));
	wire w44144;
	repeater #(2, 1'b0, 0, 0) c44144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44144));
	wire w49144;
	repeater #(2, 1'b0, 0, 0) c49144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49144));
	wire w56144;
	repeater #(1, 1'b0, 0, 0) c56144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56144));
	wire w78144;
	repeater #(1, 1'b1, 0, 0) c78144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78144));
	wire w85144;
	repeater #(2, 1'b0, 0, 0) c85144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85144));
	wire w90144;
	repeater #(2, 1'b0, 0, 0) c90144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90144));
	wire w95144;
	repeater #(2, 1'b0, 0, 0) c95144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95144));
	wire w174144;
	torch #(1'b1) c174144 (.i_clk(tick), .i_in(), .o_out(w174144));
	wire w175144;

	wire w190144;
	torch #(1'b1) c190144 (.i_clk(tick), .i_in(), .o_out(w190144));
	wire w191144;

	wire w0145;
	torch #(1'b1) c0145 (.i_clk(tick), .i_in(), .o_out(w0145));
	wire w1145;

	wire w16145;
	torch #(1'b1) c16145 (.i_clk(tick), .i_in(), .o_out(w16145));
	wire w17145;

	wire w67145;

	wire w175145;

	wire w177145;

	wire w191145;

	wire w193145;

	wire w1146;

	wire w3146;

	wire w17146;

	wire w19146;

	wire w38146;

	wire w39146;

	wire w68146;

	wire w95146;

	wire w96146;

	wire w42147;
	repeater #(2, 1'b1, 0, 0) c42147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42147));
	wire w43147;
	repeater #(2, 1'b1, 0, 0) c43147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43147));
	wire w45147;

	wire w59147;
	repeater #(1, 1'b0, 0, 0) c59147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59147));
	wire w60147;

	wire w68147;
	repeater #(1, 1'b0, 0, 0) c68147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68147));
	wire w74147;

	wire w75147;
	repeater #(1, 1'b1, 0, 0) c75147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75147));
	wire w89147;

	wire w91147;
	repeater #(2, 1'b0, 0, 0) c91147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91147));
	wire w92147;
	repeater #(2, 1'b0, 0, 0) c92147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92147));
	wire w177147;

	wire w178147;

	wire w179147;

	wire w193147;

	wire w194147;

	wire w195147;

	wire w3148;

	wire w4148;

	wire w5148;

	wire w19148;

	wire w20148;

	wire w21148;

	wire w43148;

	wire w45148;
	repeater #(1, 1'b1, 0, 0) c45148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45148));
	wire w56148;

	wire w57148;

	wire w77148;

	wire w78148;

	wire w89148;
	repeater #(1, 1'b0, 0, 0) c89148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89148));
	wire w91148;

	wire w105148;
	torch #(1'b1) c105148 (.i_clk(tick), .i_in(), .o_out(w105148));
	wire w109148;
	torch #(1'b1) c109148 (.i_clk(tick), .i_in(), .o_out(w109148));
	wire w113148;
	torch #(1'b1) c113148 (.i_clk(tick), .i_in(), .o_out(w113148));
	wire w117148;
	torch #(1'b0) c117148 (.i_clk(tick), .i_in(), .o_out(w117148));
	wire w121148;
	torch #(1'b1) c121148 (.i_clk(tick), .i_in(), .o_out(w121148));
	wire w125148;
	torch #(1'b1) c125148 (.i_clk(tick), .i_in(), .o_out(w125148));
	wire w129148;
	torch #(1'b1) c129148 (.i_clk(tick), .i_in(), .o_out(w129148));
	wire w179148;

	wire w188148;

	wire w189148;

	wire w195148;

	wire w5149;

	wire w14149;

	wire w15149;

	wire w21149;

	wire w39149;

	wire w43149;

	wire w67149;

	wire w68149;

	wire w91149;

	wire w95149;

	wire w106149;
	repeater #(1, 1'b0, 0, 0) c106149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106149));
	wire w110149;
	repeater #(1, 1'b0, 0, 0) c110149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110149));
	wire w114149;
	repeater #(1, 1'b0, 0, 0) c114149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114149));
	wire w118149;
	repeater #(1, 1'b1, 0, 0) c118149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118149));
	wire w122149;
	repeater #(1, 1'b0, 0, 0) c122149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122149));
	wire w126149;
	repeater #(1, 1'b0, 0, 0) c126149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126149));
	wire w130149;
	repeater #(1, 1'b0, 0, 0) c130149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130149));
	wire w39150;

	wire w41150;
	repeater #(1, 1'b0, 0, 0) c41150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41150));
	wire w46150;

	wire w50150;

	wire w56150;
	repeater #(1, 1'b0, 0, 0) c56150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56150));
	wire w64150;

	wire w65150;
	repeater #(1, 1'b0, 0, 0) c65150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65150));
	wire w78150;
	repeater #(1, 1'b1, 0, 0) c78150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78150));
	wire w84150;

	wire w88150;

	wire w93150;
	repeater #(1, 1'b0, 0, 0) c93150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93150));
	wire w95150;

	wire w177150;
	repeater #(1, 1'b0, 0, 0) c177150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177150));
	wire w179150;
	torch #(1'b0) c179150 (.i_clk(tick), .i_in(), .o_out(w179150));
	wire w185150;
	torch #(1'b0) c185150 (.i_clk(tick), .i_in(), .o_out(w185150));
	wire w193150;
	repeater #(1, 1'b0, 0, 0) c193150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193150));
	wire w195150;
	torch #(1'b0) c195150 (.i_clk(tick), .i_in(), .o_out(w195150));
	wire w201150;
	torch #(1'b0) c201150 (.i_clk(tick), .i_in(), .o_out(w201150));
	wire w3151;
	repeater #(1, 1'b0, 0, 0) c3151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3151));
	wire w5151;
	torch #(1'b0) c5151 (.i_clk(tick), .i_in(), .o_out(w5151));
	wire w11151;
	torch #(1'b0) c11151 (.i_clk(tick), .i_in(), .o_out(w11151));
	wire w19151;
	repeater #(1, 1'b0, 0, 0) c19151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19151));
	wire w21151;
	torch #(1'b0) c21151 (.i_clk(tick), .i_in(), .o_out(w21151));
	wire w27151;
	torch #(1'b0) c27151 (.i_clk(tick), .i_in(), .o_out(w27151));
	wire w46151;

	wire w48151;
	repeater #(1, 1'b1, 0, 0) c48151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48151));
	wire w49151;

	wire w56151;

	wire w73151;

	wire w78151;

	wire w85151;

	wire w86151;
	repeater #(1, 1'b0, 0, 0) c86151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86151));
	wire w88151;

	wire w104151;

	wire w106151;
	repeater #(1, 1'b0, 0, 0) c106151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106151));
	wire w108151;

	wire w110151;
	repeater #(1, 1'b0, 0, 0) c110151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110151));
	wire w112151;

	wire w114151;
	repeater #(1, 1'b0, 0, 0) c114151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114151));
	wire w116151;

	wire w118151;
	repeater #(1, 1'b1, 0, 0) c118151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118151));
	wire w120151;

	wire w122151;
	repeater #(1, 1'b0, 0, 0) c122151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122151));
	wire w124151;

	wire w126151;
	repeater #(1, 1'b0, 0, 0) c126151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126151));
	wire w128151;

	wire w130151;
	repeater #(1, 1'b0, 0, 0) c130151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130151));
	wire w42152;

	wire w57152;

	wire w61152;
	repeater #(1, 1'b0, 0, 0) c61152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61152));
	wire w74152;
	repeater #(2, 1'b1, 0, 0) c74152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74152));
	wire w77152;

	wire w92152;

	wire w181152;
	repeater #(1, 1'b1, 0, 0) c181152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181152));
	wire w197152;
	repeater #(1, 1'b1, 0, 0) c197152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197152));
	wire w7153;
	repeater #(1, 1'b1, 0, 0) c7153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7153));
	wire w23153;
	repeater #(1, 1'b1, 0, 0) c23153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23153));
	wire w39153;

	wire w40153;
	repeater #(1, 1'b0, 0, 0) c40153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40153));
	wire w47153;
	repeater #(2, 1'b1, 0, 0) c47153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47153));
	wire w60153;
	assign outputs[16] = ();
	wire w87153;
	repeater #(2, 1'b0, 0, 0) c87153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87153));
	wire w94153;
	repeater #(1, 1'b0, 0, 0) c94153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94153));
	wire w95153;

	wire w178154;
	torch #(1'b1) c178154 (.i_clk(tick), .i_in(), .o_out(w178154));
	wire w194154;
	torch #(1'b1) c194154 (.i_clk(tick), .i_in(), .o_out(w194154));
	wire w4155;
	torch #(1'b1) c4155 (.i_clk(tick), .i_in(), .o_out(w4155));
	wire w20155;
	torch #(1'b1) c20155 (.i_clk(tick), .i_in(), .o_out(w20155));
	wire w112155;
	torch #(1'b1) c112155 (.i_clk(tick), .i_in(), .o_out(w112155));
	wire w116155;
	torch #(1'b1) c116155 (.i_clk(tick), .i_in(), .o_out(w116155));
	wire w120155;
	torch #(1'b1) c120155 (.i_clk(tick), .i_in(), .o_out(w120155));
	wire w124155;
	torch #(1'b1) c124155 (.i_clk(tick), .i_in(), .o_out(w124155));
	wire w186156;
	torch #(1'b1) c186156 (.i_clk(tick), .i_in(), .o_out(w186156));
	wire w202156;
	torch #(1'b1) c202156 (.i_clk(tick), .i_in(), .o_out(w202156));
	wire w12157;
	torch #(1'b1) c12157 (.i_clk(tick), .i_in(), .o_out(w12157));
	wire w28157;
	torch #(1'b1) c28157 (.i_clk(tick), .i_in(), .o_out(w28157));
	wire w177157;
	repeater #(1, 1'b0, 0, 0) c177157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177157));
	wire w193157;
	repeater #(1, 1'b0, 0, 0) c193157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193157));
	wire w3158;
	repeater #(1, 1'b0, 0, 0) c3158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3158));
	wire w19158;
	repeater #(1, 1'b0, 0, 0) c19158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19158));
	wire w187158;
	repeater #(1, 1'b0, 0, 0) c187158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187158));
	wire w203158;
	repeater #(1, 1'b0, 0, 0) c203158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203158));
	wire w13159;
	repeater #(1, 1'b0, 0, 0) c13159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13159));
	wire w29159;
	repeater #(1, 1'b0, 0, 0) c29159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29159));
	wire w105164;
	torch #(1'b1) c105164 (.i_clk(tick), .i_in(), .o_out(w105164));
	wire w109164;
	torch #(1'b1) c109164 (.i_clk(tick), .i_in(), .o_out(w109164));
	wire w113164;
	torch #(1'b1) c113164 (.i_clk(tick), .i_in(), .o_out(w113164));
	wire w117164;
	torch #(1'b1) c117164 (.i_clk(tick), .i_in(), .o_out(w117164));
	wire w121164;
	torch #(1'b1) c121164 (.i_clk(tick), .i_in(), .o_out(w121164));
	wire w125164;
	torch #(1'b1) c125164 (.i_clk(tick), .i_in(), .o_out(w125164));
	wire w129164;
	torch #(1'b1) c129164 (.i_clk(tick), .i_in(), .o_out(w129164));
	wire w106165;
	repeater #(1, 1'b0, 0, 0) c106165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106165));
	wire w110165;
	repeater #(1, 1'b0, 0, 0) c110165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110165));
	wire w114165;
	repeater #(1, 1'b0, 0, 0) c114165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114165));
	wire w118165;
	repeater #(1, 1'b1, 0, 0) c118165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118165));
	wire w122165;
	repeater #(1, 1'b0, 0, 0) c122165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122165));
	wire w126165;
	repeater #(1, 1'b0, 0, 0) c126165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126165));
	wire w130165;
	repeater #(1, 1'b0, 0, 0) c130165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130165));
	wire w104167;

	wire w106167;
	repeater #(1, 1'b0, 0, 0) c106167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106167));
	wire w108167;

	wire w110167;
	repeater #(1, 1'b0, 0, 0) c110167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110167));
	wire w112167;

	wire w114167;
	repeater #(1, 1'b0, 0, 0) c114167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114167));
	wire w116167;

	wire w118167;
	repeater #(1, 1'b1, 0, 0) c118167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118167));
	wire w120167;

	wire w122167;
	repeater #(1, 1'b0, 0, 0) c122167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122167));
	wire w124167;

	wire w126167;
	repeater #(1, 1'b0, 0, 0) c126167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126167));
	wire w128167;

	wire w130167;
	repeater #(1, 1'b0, 0, 0) c130167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130167));
	wire w112171;
	torch #(1'b1) c112171 (.i_clk(tick), .i_in(), .o_out(w112171));
	wire w116171;
	torch #(1'b1) c116171 (.i_clk(tick), .i_in(), .o_out(w116171));
	wire w120171;
	torch #(1'b1) c120171 (.i_clk(tick), .i_in(), .o_out(w120171));
	wire w124171;
	torch #(1'b1) c124171 (.i_clk(tick), .i_in(), .o_out(w124171));
	wire w66175;

	wire w67175;
	repeater #(1, 1'b0, 0, 0) c67175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67175));
	wire w68176;
	repeater #(1, 1'b0, 0, 0) c68176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68176));
	wire w71176;
	repeater #(2, 1'b0, 0, 0) c71176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71176));
	wire w63177;
	repeater #(1, 1'b0, 0, 0) c63177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63177));
	wire w76177;
	repeater #(2, 1'b0, 0, 0) c76177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76177));
	wire w62178;
	assign outputs[17] = ();
	wire w65178;

	wire w74178;

	wire w65179;

	wire w74179;

	wire w63180;
	repeater #(1, 1'b0, 0, 0) c63180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63180));
	wire w76180;
	repeater #(1, 1'b0, 0, 0) c76180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76180));
	wire w105180;
	torch #(1'b1) c105180 (.i_clk(tick), .i_in(), .o_out(w105180));
	wire w109180;
	torch #(1'b1) c109180 (.i_clk(tick), .i_in(), .o_out(w109180));
	wire w113180;
	torch #(1'b1) c113180 (.i_clk(tick), .i_in(), .o_out(w113180));
	wire w117180;
	torch #(1'b0) c117180 (.i_clk(tick), .i_in(), .o_out(w117180));
	wire w121180;
	torch #(1'b1) c121180 (.i_clk(tick), .i_in(), .o_out(w121180));
	wire w125180;
	torch #(1'b1) c125180 (.i_clk(tick), .i_in(), .o_out(w125180));
	wire w129180;
	torch #(1'b1) c129180 (.i_clk(tick), .i_in(), .o_out(w129180));
	wire w106181;
	repeater #(1, 1'b0, 0, 0) c106181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106181));
	wire w110181;
	repeater #(1, 1'b0, 0, 0) c110181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110181));
	wire w114181;
	repeater #(1, 1'b0, 0, 0) c114181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114181));
	wire w118181;
	repeater #(1, 1'b1, 0, 0) c118181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118181));
	wire w122181;
	repeater #(1, 1'b0, 0, 0) c122181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122181));
	wire w126181;
	repeater #(1, 1'b0, 0, 0) c126181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126181));
	wire w130181;
	repeater #(1, 1'b0, 0, 0) c130181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130181));
	wire w104183;

	wire w106183;
	repeater #(1, 1'b0, 0, 0) c106183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106183));
	wire w108183;

	wire w110183;
	repeater #(1, 1'b0, 0, 0) c110183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110183));
	wire w112183;

	wire w114183;
	repeater #(1, 1'b0, 0, 0) c114183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114183));
	wire w116183;

	wire w118183;
	repeater #(1, 1'b1, 0, 0) c118183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118183));
	wire w120183;

	wire w122183;
	repeater #(1, 1'b0, 0, 0) c122183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122183));
	wire w124183;

	wire w126183;
	repeater #(1, 1'b0, 0, 0) c126183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126183));
	wire w128183;

	wire w130183;
	repeater #(1, 1'b0, 0, 0) c130183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130183));
	wire w112187;
	torch #(1'b1) c112187 (.i_clk(tick), .i_in(), .o_out(w112187));
	wire w116187;
	torch #(1'b1) c116187 (.i_clk(tick), .i_in(), .o_out(w116187));
	wire w120187;
	torch #(1'b1) c120187 (.i_clk(tick), .i_in(), .o_out(w120187));
	wire w124187;
	torch #(1'b1) c124187 (.i_clk(tick), .i_in(), .o_out(w124187));
	wire w105196;
	torch #(1'b1) c105196 (.i_clk(tick), .i_in(), .o_out(w105196));
	wire w109196;
	torch #(1'b1) c109196 (.i_clk(tick), .i_in(), .o_out(w109196));
	wire w113196;
	torch #(1'b1) c113196 (.i_clk(tick), .i_in(), .o_out(w113196));
	wire w117196;
	torch #(1'b1) c117196 (.i_clk(tick), .i_in(), .o_out(w117196));
	wire w121196;
	torch #(1'b1) c121196 (.i_clk(tick), .i_in(), .o_out(w121196));
	wire w125196;
	torch #(1'b1) c125196 (.i_clk(tick), .i_in(), .o_out(w125196));
	wire w129196;
	torch #(1'b1) c129196 (.i_clk(tick), .i_in(), .o_out(w129196));
	wire w106197;
	repeater #(1, 1'b0, 0, 0) c106197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106197));
	wire w110197;
	repeater #(1, 1'b0, 0, 0) c110197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110197));
	wire w114197;
	repeater #(1, 1'b0, 0, 0) c114197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114197));
	wire w118197;
	repeater #(1, 1'b1, 0, 0) c118197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118197));
	wire w122197;
	repeater #(1, 1'b0, 0, 0) c122197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122197));
	wire w126197;
	repeater #(1, 1'b0, 0, 0) c126197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126197));
	wire w130197;
	repeater #(1, 1'b0, 0, 0) c130197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130197));
	wire w104199;

	wire w106199;
	repeater #(1, 1'b0, 0, 0) c106199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106199));
	wire w108199;

	wire w110199;
	repeater #(1, 1'b0, 0, 0) c110199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110199));
	wire w112199;

	wire w114199;
	repeater #(1, 1'b0, 0, 0) c114199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114199));
	wire w116199;

	wire w118199;
	repeater #(1, 1'b1, 0, 0) c118199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118199));
	wire w120199;

	wire w122199;
	repeater #(1, 1'b0, 0, 0) c122199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122199));
	wire w124199;

	wire w126199;
	repeater #(1, 1'b0, 0, 0) c126199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126199));
	wire w128199;

	wire w130199;
	repeater #(1, 1'b0, 0, 0) c130199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130199));
	wire w1051105;
	torch #(1'b1) c1051105 (.i_clk(tick), .i_in(), .o_out(w1051105));
	wire w1091105;
	torch #(1'b1) c1091105 (.i_clk(tick), .i_in(), .o_out(w1091105));
	wire w1131105;
	torch #(1'b1) c1131105 (.i_clk(tick), .i_in(), .o_out(w1131105));
	wire w1171105;
	torch #(1'b0) c1171105 (.i_clk(tick), .i_in(), .o_out(w1171105));
	wire w1211105;
	torch #(1'b1) c1211105 (.i_clk(tick), .i_in(), .o_out(w1211105));
	wire w1251105;
	torch #(1'b1) c1251105 (.i_clk(tick), .i_in(), .o_out(w1251105));
	wire w1291105;
	torch #(1'b1) c1291105 (.i_clk(tick), .i_in(), .o_out(w1291105));
	wire w1061117;
	repeater #(1, 1'b0, 0, 0) c1061117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061117));
	wire w1101117;
	repeater #(1, 1'b0, 0, 0) c1101117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101117));
	wire w1141117;
	repeater #(1, 1'b0, 0, 0) c1141117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1141117));
	wire w1181117;
	repeater #(1, 1'b1, 0, 0) c1181117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1181117));
	wire w1221117;
	repeater #(1, 1'b0, 0, 0) c1221117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221117));
	wire w1261117;
	repeater #(1, 1'b0, 0, 0) c1261117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1261117));
	wire w1301117;
	repeater #(1, 1'b0, 0, 0) c1301117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1301117));
	wire w1051118;
	repeater #(1, 1'b1, 0, 0) c1051118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1051118));
	wire w1091118;
	repeater #(1, 1'b1, 0, 0) c1091118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1091118));
	wire w1131118;
	repeater #(1, 1'b0, 0, 0) c1131118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1131118));
	wire w1171118;
	repeater #(1, 1'b1, 0, 0) c1171118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1171118));
	wire w1211118;
	repeater #(1, 1'b0, 0, 0) c1211118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1211118));
	wire w1251118;
	repeater #(1, 1'b1, 0, 0) c1251118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1251118));
	wire w1291118;
	repeater #(1, 1'b1, 0, 0) c1291118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1291118));
	wire w1331118;
	torch #(1'b0) c1331118 (.i_clk(tick), .i_in(), .o_out(w1331118));
	wire w1041122;
	torch #(1'b0) c1041122 (.i_clk(tick), .i_in(), .o_out(w1041122));
	wire w1081122;
	torch #(1'b0) c1081122 (.i_clk(tick), .i_in(), .o_out(w1081122));
	wire w1121122;
	torch #(1'b0) c1121122 (.i_clk(tick), .i_in(), .o_out(w1121122));
	wire w1161122;
	torch #(1'b0) c1161122 (.i_clk(tick), .i_in(), .o_out(w1161122));
	wire w1201122;
	torch #(1'b0) c1201122 (.i_clk(tick), .i_in(), .o_out(w1201122));
	wire w1241122;
	torch #(1'b0) c1241122 (.i_clk(tick), .i_in(), .o_out(w1241122));
	wire w1281122;
	torch #(1'b0) c1281122 (.i_clk(tick), .i_in(), .o_out(w1281122));
	wire w1351124;
	torch #(1'b1) c1351124 (.i_clk(tick), .i_in(), .o_out(w1351124));
	wire w89016;
	torch #(1'b1) c89016 (.i_clk(tick), .i_in(), .o_out(w89016));
	wire w93016;
	torch #(1'b1) c93016 (.i_clk(tick), .i_in(), .o_out(w93016));
	wire w97016;
	torch #(1'b1) c97016 (.i_clk(tick), .i_in(), .o_out(w97016));
	wire w101016;
	torch #(1'b0) c101016 (.i_clk(tick), .i_in(), .o_out(w101016));
	wire w105016;
	torch #(1'b1) c105016 (.i_clk(tick), .i_in(), .o_out(w105016));
	wire w109016;
	torch #(1'b1) c109016 (.i_clk(tick), .i_in(), .o_out(w109016));
	wire w113016;
	torch #(1'b1) c113016 (.i_clk(tick), .i_in(), .o_out(w113016));
	wire w205020;

	wire w31021;

	wire w65021;

	wire w99021;

	wire w204021;
	repeater #(1, 1'b1, 0, 0) c204021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204021));
	wire w30022;
	repeater #(1, 1'b1, 0, 0) c30022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30022));
	wire w64022;
	repeater #(1, 1'b1, 0, 0) c64022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64022));
	wire w98022;
	repeater #(1, 1'b1, 0, 0) c98022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98022));
	wire w203022;

	wire w29023;

	wire w63023;

	wire w97023;

	wire w202023;
	repeater #(1, 1'b1, 0, 0) c202023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202023));
	wire w28024;
	repeater #(1, 1'b1, 0, 0) c28024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28024));
	wire w62024;
	repeater #(1, 1'b1, 0, 0) c62024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62024));
	wire w96024;
	repeater #(1, 1'b1, 0, 0) c96024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96024));
	wire w201024;

	wire w27025;

	wire w61025;

	wire w95025;

	wire w200025;
	repeater #(1, 1'b1, 0, 0) c200025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200025));
	wire w26026;
	repeater #(1, 1'b1, 0, 0) c26026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26026));
	wire w60026;
	repeater #(1, 1'b1, 0, 0) c60026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60026));
	wire w94026;
	repeater #(1, 1'b1, 0, 0) c94026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94026));
	wire w199026;

	wire w25027;

	wire w59027;

	wire w93027;

	wire w198027;
	repeater #(1, 1'b1, 0, 0) c198027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198027));
	wire w24028;
	repeater #(1, 1'b1, 0, 0) c24028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24028));
	wire w58028;
	repeater #(1, 1'b1, 0, 0) c58028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58028));
	wire w92028;
	repeater #(1, 1'b1, 0, 0) c92028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92028));
	wire w197028;

	wire w23029;

	wire w57029;

	wire w91029;

	wire w196029;
	repeater #(1, 1'b1, 0, 0) c196029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196029));
	wire w22030;
	repeater #(1, 1'b1, 0, 0) c22030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22030));
	wire w56030;
	repeater #(1, 1'b1, 0, 0) c56030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56030));
	wire w90030;
	repeater #(1, 1'b1, 0, 0) c90030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90030));
	wire w195030;

	wire w21031;

	wire w55031;

	wire w89031;

	wire w194031;
	repeater #(1, 1'b1, 0, 0) c194031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194031));
	wire w20032;
	repeater #(1, 1'b1, 0, 0) c20032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20032));
	wire w54032;
	repeater #(1, 1'b1, 0, 0) c54032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54032));
	wire w88032;
	repeater #(1, 1'b1, 0, 0) c88032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88032));
	wire w193032;

	wire w19033;

	wire w53033;

	wire w87033;

	wire w192033;
	repeater #(1, 1'b0, 0, 0) c192033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192033));
	wire w18034;
	repeater #(1, 1'b0, 0, 0) c18034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18034));
	wire w52034;
	repeater #(1, 1'b0, 0, 0) c52034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52034));
	wire w86034;
	repeater #(1, 1'b0, 0, 0) c86034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86034));
	wire w191034;

	wire w17035;

	wire w51035;

	wire w85035;

	wire w190035;
	repeater #(1, 1'b0, 0, 0) c190035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190035));
	wire w16036;
	repeater #(1, 1'b0, 0, 0) c16036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16036));
	wire w50036;
	repeater #(1, 1'b0, 0, 0) c50036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50036));
	wire w84036;
	repeater #(1, 1'b0, 0, 0) c84036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84036));
	wire w189036;

	wire w15037;

	wire w49037;

	wire w83037;

	wire w188037;
	repeater #(1, 1'b1, 0, 0) c188037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188037));
	wire w14038;
	repeater #(1, 1'b1, 0, 0) c14038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14038));
	wire w48038;
	repeater #(1, 1'b1, 0, 0) c48038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48038));
	wire w82038;
	repeater #(1, 1'b1, 0, 0) c82038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82038));
	wire w187038;

	wire w13039;

	wire w47039;

	wire w81039;

	wire w186039;
	repeater #(1, 1'b1, 0, 0) c186039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186039));
	wire w12040;
	repeater #(1, 1'b1, 0, 0) c12040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12040));
	wire w46040;
	repeater #(1, 1'b1, 0, 0) c46040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46040));
	wire w80040;
	repeater #(1, 1'b1, 0, 0) c80040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80040));
	wire w185040;

	wire w11041;

	wire w45041;

	wire w79041;

	wire w184041;
	repeater #(1, 1'b1, 0, 0) c184041 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184041));
	wire w10042;
	repeater #(1, 1'b1, 0, 0) c10042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10042));
	wire w44042;
	repeater #(1, 1'b1, 0, 0) c44042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44042));
	wire w78042;
	repeater #(1, 1'b1, 0, 0) c78042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78042));
	wire w183042;

	wire w9043;

	wire w43043;

	wire w77043;

	wire w182043;
	repeater #(1, 1'b1, 0, 0) c182043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182043));
	wire w8044;
	repeater #(1, 1'b1, 0, 0) c8044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8044));
	wire w42044;
	repeater #(1, 1'b1, 0, 0) c42044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42044));
	wire w76044;
	repeater #(1, 1'b1, 0, 0) c76044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76044));
	wire w181044;

	wire w7045;

	wire w41045;

	wire w75045;

	wire w180045;
	repeater #(1, 1'b1, 0, 0) c180045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180045));
	wire w6046;
	repeater #(1, 1'b1, 0, 0) c6046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6046));
	wire w40046;
	repeater #(1, 1'b1, 0, 0) c40046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40046));
	wire w74046;
	repeater #(1, 1'b1, 0, 0) c74046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74046));
	wire w179046;

	wire w5047;

	wire w39047;

	wire w73047;

	wire w178047;
	repeater #(1, 1'b1, 0, 0) c178047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178047));
	wire w4048;
	repeater #(1, 1'b1, 0, 0) c4048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4048));
	wire w38048;
	repeater #(1, 1'b1, 0, 0) c38048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38048));
	wire w72048;
	repeater #(1, 1'b1, 0, 0) c72048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72048));
	wire w176052;
	repeater #(2, 1'b1, 0, 0) c176052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176052));
	wire w2053;
	repeater #(2, 1'b1, 0, 0) c2053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2053));
	wire w88054;
	repeater #(1, 1'b1, 0, 0) c88054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88054));
	wire w92054;
	repeater #(1, 1'b1, 0, 0) c92054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92054));
	wire w96054;
	repeater #(1, 1'b1, 0, 0) c96054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96054));
	wire w100054;
	repeater #(1, 1'b0, 0, 0) c100054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100054));
	wire w104054;
	repeater #(1, 1'b1, 0, 0) c104054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104054));
	wire w108054;
	repeater #(1, 1'b1, 0, 0) c108054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108054));
	wire w112054;
	repeater #(1, 1'b1, 0, 0) c112054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112054));
	wire w162054;
	repeater #(1, 1'b1, 0, 0) c162054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162054));
	wire w168054;
	torch #(1'b1) c168054 (.i_clk(tick), .i_in(), .o_out(w168054));
	wire w178054;
	repeater #(1, 1'b1, 0, 0) c178054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178054));
	wire w184054;
	torch #(1'b1) c184054 (.i_clk(tick), .i_in(), .o_out(w184054));
	wire w196054;
	repeater #(1, 1'b1, 0, 0) c196054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196054));
	wire w202054;
	torch #(1'b1) c202054 (.i_clk(tick), .i_in(), .o_out(w202054));
	wire w4055;
	repeater #(1, 1'b1, 0, 0) c4055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4055));
	wire w10055;
	torch #(1'b1) c10055 (.i_clk(tick), .i_in(), .o_out(w10055));
	wire w88055;
	repeater #(1, 1'b1, 0, 0) c88055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88055));
	wire w90055;
	repeater #(1, 1'b0, 0, 0) c90055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90055));
	wire w92055;
	repeater #(1, 1'b1, 0, 0) c92055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92055));
	wire w94055;
	repeater #(1, 1'b0, 0, 0) c94055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94055));
	wire w96055;
	repeater #(1, 1'b1, 0, 0) c96055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96055));
	wire w98055;
	repeater #(1, 1'b0, 0, 0) c98055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98055));
	wire w100055;
	repeater #(1, 1'b0, 0, 0) c100055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100055));
	wire w102055;
	repeater #(1, 1'b0, 0, 0) c102055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102055));
	wire w104055;
	repeater #(1, 1'b1, 0, 0) c104055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104055));
	wire w106055;
	repeater #(1, 1'b0, 0, 0) c106055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106055));
	wire w108055;
	repeater #(1, 1'b1, 0, 0) c108055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108055));
	wire w110055;
	repeater #(1, 1'b0, 0, 0) c110055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110055));
	wire w112055;
	repeater #(1, 1'b1, 0, 0) c112055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112055));
	wire w114055;
	repeater #(1, 1'b0, 0, 0) c114055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114055));
	wire w89056;
	torch #(1'b0) c89056 (.i_clk(tick), .i_in(), .o_out(w89056));
	wire w93056;
	torch #(1'b0) c93056 (.i_clk(tick), .i_in(), .o_out(w93056));
	wire w97056;
	torch #(1'b0) c97056 (.i_clk(tick), .i_in(), .o_out(w97056));
	wire w101056;
	torch #(1'b0) c101056 (.i_clk(tick), .i_in(), .o_out(w101056));
	wire w105056;
	torch #(1'b0) c105056 (.i_clk(tick), .i_in(), .o_out(w105056));
	wire w109056;
	torch #(1'b0) c109056 (.i_clk(tick), .i_in(), .o_out(w109056));
	wire w113056;
	torch #(1'b0) c113056 (.i_clk(tick), .i_in(), .o_out(w113056));
	wire w169057;
	repeater #(1, 1'b1, 0, 0) c169057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169057));
	wire w185057;
	repeater #(1, 1'b1, 0, 0) c185057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185057));
	wire w203057;
	repeater #(1, 1'b1, 0, 0) c203057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203057));
	wire w11058;
	repeater #(1, 1'b1, 0, 0) c11058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11058));
	wire w162058;
	repeater #(1, 1'b1, 0, 0) c162058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162058));
	wire w178058;
	repeater #(1, 1'b1, 0, 0) c178058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178058));
	wire w196058;
	repeater #(1, 1'b1, 0, 0) c196058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196058));
	wire w4059;
	repeater #(1, 1'b1, 0, 0) c4059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4059));
	wire w29059;
	repeater #(1, 1'b0, 0, 0) c29059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29059));
	wire w33059;
	repeater #(1, 1'b0, 0, 0) c33059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33059));
	wire w37059;
	repeater #(1, 1'b0, 0, 0) c37059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37059));
	wire w41059;
	repeater #(1, 1'b0, 0, 0) c41059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41059));
	wire w61059;
	repeater #(1, 1'b1, 0, 0) c61059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61059));
	wire w65059;
	repeater #(1, 1'b1, 0, 0) c65059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65059));
	wire w69059;
	repeater #(1, 1'b1, 0, 0) c69059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69059));
	wire w73059;
	repeater #(1, 1'b1, 0, 0) c73059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73059));
	wire w167059;

	wire w183059;

	wire w201059;

	wire w9060;

	wire w175060;

	wire w1061;

	wire w161061;

	wire w162061;

	wire w172061;

	wire w177061;

	wire w178061;

	wire w195061;

	wire w196061;

	wire w206061;

	wire w3062;

	wire w4062;

	wire w27062;
	torch #(1'b1) c27062 (.i_clk(tick), .i_in(), .o_out(w27062));
	wire w31062;
	torch #(1'b1) c31062 (.i_clk(tick), .i_in(), .o_out(w31062));
	wire w35062;
	torch #(1'b0) c35062 (.i_clk(tick), .i_in(), .o_out(w35062));
	wire w39062;
	torch #(1'b1) c39062 (.i_clk(tick), .i_in(), .o_out(w39062));
	wire w63062;
	torch #(1'b0) c63062 (.i_clk(tick), .i_in(), .o_out(w63062));
	wire w67062;
	torch #(1'b1) c67062 (.i_clk(tick), .i_in(), .o_out(w67062));
	wire w71062;
	torch #(1'b0) c71062 (.i_clk(tick), .i_in(), .o_out(w71062));
	wire w75062;
	torch #(1'b0) c75062 (.i_clk(tick), .i_in(), .o_out(w75062));
	wire w96063;
	torch #(1'b1) c96063 (.i_clk(tick), .i_in(), .o_out(w96063));
	wire w100063;
	torch #(1'b1) c100063 (.i_clk(tick), .i_in(), .o_out(w100063));
	wire w104063;
	torch #(1'b1) c104063 (.i_clk(tick), .i_in(), .o_out(w104063));
	wire w108063;
	torch #(1'b1) c108063 (.i_clk(tick), .i_in(), .o_out(w108063));
	wire w170063;

	wire w204063;

	wire w160064;

	wire w161064;

	wire w176064;

	wire w177064;

	wire w194064;

	wire w195064;

	wire w2065;

	wire w3065;

	wire w162065;

	wire w166065;

	wire w170065;

	wire w196065;

	wire w200065;

	wire w204065;

	wire w90066;

	wire w94066;

	wire w98066;

	wire w102066;

	wire w106066;

	wire w110066;

	wire w114066;

	wire w186068;

	wire w12069;

	wire w159069;

	wire w160069;

	wire w163069;

	wire w164069;

	wire w167069;

	wire w168069;

	wire w171069;

	wire w172069;

	wire w175069;

	wire w176069;

	wire w179069;

	wire w180069;

	wire w183069;

	wire w184069;

	wire w193069;

	wire w194069;

	wire w197069;

	wire w198069;

	wire w201069;

	wire w202069;

	wire w205069;

	wire w206069;

	wire w1070;

	wire w2070;

	wire w5070;

	wire w6070;

	wire w9070;

	wire w10070;

	wire w157070;

	wire w191070;

	wire w172073;
	repeater #(1, 1'b1, 0, 0) c172073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172073));
	wire w176073;
	repeater #(1, 1'b1, 0, 0) c176073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176073));
	wire w180073;
	repeater #(1, 1'b1, 0, 0) c180073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180073));
	wire w206073;
	repeater #(1, 1'b1, 0, 0) c206073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206073));
	wire w2074;
	repeater #(1, 1'b1, 0, 0) c2074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2074));
	wire w6074;
	repeater #(1, 1'b1, 0, 0) c6074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6074));
	wire w91075;
	torch #(1'b0) c91075 (.i_clk(tick), .i_in(), .o_out(w91075));
	wire w95075;
	torch #(1'b0) c95075 (.i_clk(tick), .i_in(), .o_out(w95075));
	wire w99075;
	torch #(1'b0) c99075 (.i_clk(tick), .i_in(), .o_out(w99075));
	wire w103075;
	torch #(1'b0) c103075 (.i_clk(tick), .i_in(), .o_out(w103075));
	wire w107075;
	torch #(1'b0) c107075 (.i_clk(tick), .i_in(), .o_out(w107075));
	wire w111075;
	torch #(1'b0) c111075 (.i_clk(tick), .i_in(), .o_out(w111075));
	wire w115075;
	torch #(1'b0) c115075 (.i_clk(tick), .i_in(), .o_out(w115075));
	wire w158076;

	wire w162076;

	wire w178076;

	wire w182076;

	wire w192076;

	wire w196076;

	wire w4077;

	wire w8077;

	wire w90077;
	torch #(1'b0) c90077 (.i_clk(tick), .i_in(), .o_out(w90077));
	wire w94077;
	torch #(1'b0) c94077 (.i_clk(tick), .i_in(), .o_out(w94077));
	wire w98077;
	torch #(1'b0) c98077 (.i_clk(tick), .i_in(), .o_out(w98077));
	wire w102077;
	torch #(1'b1) c102077 (.i_clk(tick), .i_in(), .o_out(w102077));
	wire w106077;
	torch #(1'b0) c106077 (.i_clk(tick), .i_in(), .o_out(w106077));
	wire w110077;
	torch #(1'b0) c110077 (.i_clk(tick), .i_in(), .o_out(w110077));
	wire w114077;
	torch #(1'b0) c114077 (.i_clk(tick), .i_in(), .o_out(w114077));
	wire w160077;
	repeater #(1, 1'b1, 0, 0) c160077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160077));
	wire w176077;
	repeater #(1, 1'b1, 0, 0) c176077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176077));
	wire w194077;
	repeater #(1, 1'b1, 0, 0) c194077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194077));
	wire w2078;
	repeater #(1, 1'b1, 0, 0) c2078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2078));
	wire w154078;

	wire w167078;
	repeater #(1, 1'b0, 0, 0) c167078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167078));
	wire w188078;

	wire w201078;
	repeater #(1, 1'b1, 0, 0) c201078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201078));
	wire w96079;
	torch #(1'b1) c96079 (.i_clk(tick), .i_in(), .o_out(w96079));
	wire w100079;
	torch #(1'b1) c100079 (.i_clk(tick), .i_in(), .o_out(w100079));
	wire w104079;
	torch #(1'b1) c104079 (.i_clk(tick), .i_in(), .o_out(w104079));
	wire w108079;
	torch #(1'b1) c108079 (.i_clk(tick), .i_in(), .o_out(w108079));
	wire w162079;

	wire w178079;

	wire w196079;

	wire w4080;

	wire w154080;

	wire w170080;

	wire w188080;

	wire w204080;

	wire w157081;

	wire w165081;

	wire w167081;

	wire w168081;

	wire w173081;

	wire w181081;

	wire w191081;

	wire w199081;

	wire w201081;

	wire w202081;

	wire w207081;

	wire w7082;

	wire w90082;

	wire w94082;

	wire w98082;

	wire w102082;

	wire w106082;

	wire w110082;

	wire w114082;

	wire w159083;

	wire w160083;

	wire w175083;

	wire w176083;

	wire w193083;

	wire w194083;

	wire w1084;

	wire w2084;

	wire w165085;

	wire w167085;

	wire w168085;

	wire w181085;

	wire w199085;

	wire w201085;

	wire w202085;

	wire w7086;

	wire w50086;

	wire w49087;
	repeater #(1, 1'b1, 0, 0) c49087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49087));
	wire w162087;
	torch #(1'b1) c162087 (.i_clk(tick), .i_in(), .o_out(w162087));
	wire w163087;

	wire w178087;
	torch #(1'b1) c178087 (.i_clk(tick), .i_in(), .o_out(w178087));
	wire w179087;

	wire w196087;
	torch #(1'b1) c196087 (.i_clk(tick), .i_in(), .o_out(w196087));
	wire w197087;

	wire w4088;
	torch #(1'b1) c4088 (.i_clk(tick), .i_in(), .o_out(w4088));
	wire w5088;

	wire w24088;
	repeater #(2, 1'b1, 0, 0) c24088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24088));
	wire w78088;
	repeater #(2, 1'b1, 0, 0) c78088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78088));
	wire w163088;

	wire w165088;

	wire w179088;

	wire w181088;

	wire w197088;

	wire w199088;

	wire w5089;

	wire w7089;

	wire w21089;
	repeater #(1, 1'b1, 0, 0) c21089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21089));
	wire w29089;
	repeater #(1, 1'b1, 0, 0) c29089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29089));
	wire w30089;
	repeater #(2, 1'b1, 0, 0) c30089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30089));
	wire w53089;

	wire w72089;
	repeater #(2, 1'b0, 0, 0) c72089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72089));
	wire w73089;
	repeater #(1, 1'b0, 0, 0) c73089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73089));
	wire w81089;
	repeater #(1, 1'b1, 0, 0) c81089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81089));
	wire w25090;
	repeater #(1, 1'b1, 0, 0) c25090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25090));
	wire w50090;

	wire w77090;
	repeater #(1, 1'b0, 0, 0) c77090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77090));
	wire w165090;

	wire w166090;

	wire w167090;

	wire w181090;

	wire w182090;

	wire w183090;

	wire w199090;

	wire w200090;

	wire w201090;

	wire w7091;

	wire w8091;

	wire w9091;

	wire w31091;

	wire w35091;
	repeater #(1, 1'b0, 0, 0) c35091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35091));
	wire w49091;

	wire w51091;
	repeater #(2, 1'b1, 0, 0) c51091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51091));
	wire w54091;
	repeater #(2, 1'b0, 0, 0) c54091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54091));
	wire w67091;
	repeater #(1, 1'b1, 0, 0) c67091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67091));
	wire w71091;

	wire w91091;
	torch #(1'b0) c91091 (.i_clk(tick), .i_in(), .o_out(w91091));
	wire w95091;
	torch #(1'b0) c95091 (.i_clk(tick), .i_in(), .o_out(w95091));
	wire w99091;
	torch #(1'b0) c99091 (.i_clk(tick), .i_in(), .o_out(w99091));
	wire w103091;
	torch #(1'b0) c103091 (.i_clk(tick), .i_in(), .o_out(w103091));
	wire w107091;
	torch #(1'b0) c107091 (.i_clk(tick), .i_in(), .o_out(w107091));
	wire w111091;
	torch #(1'b0) c111091 (.i_clk(tick), .i_in(), .o_out(w111091));
	wire w115091;
	torch #(1'b0) c115091 (.i_clk(tick), .i_in(), .o_out(w115091));
	wire w160091;

	wire w161091;

	wire w167091;

	wire w176091;

	wire w177091;

	wire w183091;

	wire w194091;

	wire w195091;

	wire w201091;

	wire w2092;

	wire w3092;

	wire w9092;

	wire w32092;

	wire w38092;
	repeater #(2, 1'b0, 0, 0) c38092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38092));
	wire w41092;
	repeater #(2, 1'b0, 0, 0) c41092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41092));
	wire w43092;

	wire w59092;

	wire w61092;
	repeater #(2, 1'b0, 0, 0) c61092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61092));
	wire w64092;
	repeater #(2, 1'b1, 0, 0) c64092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64092));
	wire w70092;

	wire w31093;
	repeater #(2, 1'b1, 0, 0) c31093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31093));
	wire w42093;

	wire w60093;

	wire w71093;
	repeater #(2, 1'b1, 0, 0) c71093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71093));
	wire w90093;
	torch #(1'b0) c90093 (.i_clk(tick), .i_in(), .o_out(w90093));
	wire w94093;
	torch #(1'b0) c94093 (.i_clk(tick), .i_in(), .o_out(w94093));
	wire w98093;
	torch #(1'b0) c98093 (.i_clk(tick), .i_in(), .o_out(w98093));
	wire w102093;
	torch #(1'b1) c102093 (.i_clk(tick), .i_in(), .o_out(w102093));
	wire w106093;
	torch #(1'b0) c106093 (.i_clk(tick), .i_in(), .o_out(w106093));
	wire w110093;
	torch #(1'b0) c110093 (.i_clk(tick), .i_in(), .o_out(w110093));
	wire w114093;
	torch #(1'b0) c114093 (.i_clk(tick), .i_in(), .o_out(w114093));
	wire w165093;
	repeater #(1, 1'b0, 0, 0) c165093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165093));
	wire w167093;
	torch #(1'b0) c167093 (.i_clk(tick), .i_in(), .o_out(w167093));
	wire w173093;
	torch #(1'b1) c173093 (.i_clk(tick), .i_in(), .o_out(w173093));
	wire w181093;
	repeater #(1, 1'b0, 0, 0) c181093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181093));
	wire w183093;
	torch #(1'b0) c183093 (.i_clk(tick), .i_in(), .o_out(w183093));
	wire w199093;
	repeater #(1, 1'b0, 0, 0) c199093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199093));
	wire w201093;
	torch #(1'b0) c201093 (.i_clk(tick), .i_in(), .o_out(w201093));
	wire w207093;
	torch #(1'b1) c207093 (.i_clk(tick), .i_in(), .o_out(w207093));
	wire w7094;
	repeater #(1, 1'b0, 0, 0) c7094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7094));
	wire w9094;
	torch #(1'b0) c9094 (.i_clk(tick), .i_in(), .o_out(w9094));
	wire w25094;

	wire w26094;

	wire w39094;

	wire w63094;

	wire w76094;

	wire w77094;

	wire w24095;

	wire w33095;

	wire w69095;

	wire w78095;

	wire w96095;
	torch #(1'b1) c96095 (.i_clk(tick), .i_in(), .o_out(w96095));
	wire w100095;
	torch #(1'b1) c100095 (.i_clk(tick), .i_in(), .o_out(w100095));
	wire w104095;
	torch #(1'b1) c104095 (.i_clk(tick), .i_in(), .o_out(w104095));
	wire w108095;
	torch #(1'b1) c108095 (.i_clk(tick), .i_in(), .o_out(w108095));
	wire w169095;
	repeater #(1, 1'b1, 0, 0) c169095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169095));
	wire w185095;
	repeater #(1, 1'b1, 0, 0) c185095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185095));
	wire w203095;
	repeater #(1, 1'b1, 0, 0) c203095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203095));
	wire w11096;
	repeater #(1, 1'b1, 0, 0) c11096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11096));
	wire w27096;

	wire w57096;
	assign outputs[18] = ();
	wire w75096;

	wire w166097;
	torch #(1'b1) c166097 (.i_clk(tick), .i_in(), .o_out(w166097));
	wire w182097;
	torch #(1'b1) c182097 (.i_clk(tick), .i_in(), .o_out(w182097));
	wire w200097;
	torch #(1'b1) c200097 (.i_clk(tick), .i_in(), .o_out(w200097));
	wire w8098;
	torch #(1'b1) c8098 (.i_clk(tick), .i_in(), .o_out(w8098));
	wire w90098;

	wire w94098;

	wire w98098;

	wire w102098;

	wire w106098;

	wire w110098;

	wire w114098;

	wire w174099;
	torch #(1'b1) c174099 (.i_clk(tick), .i_in(), .o_out(w174099));
	wire w00100;
	torch #(1'b1) c00100 (.i_clk(tick), .i_in(), .o_out(w00100));
	wire w1650100;
	repeater #(1, 1'b0, 0, 0) c1650100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1650100));
	wire w1810100;
	repeater #(1, 1'b0, 0, 0) c1810100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810100));
	wire w1990100;
	repeater #(1, 1'b0, 0, 0) c1990100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990100));
	wire w70101;
	repeater #(1, 1'b0, 0, 0) c70101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70101));
	wire w1750101;
	repeater #(1, 1'b0, 0, 0) c1750101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750101));
	wire w10102;
	repeater #(1, 1'b0, 0, 0) c10102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10102));
	wire w910107;
	torch #(1'b0) c910107 (.i_clk(tick), .i_in(), .o_out(w910107));
	wire w950107;
	torch #(1'b0) c950107 (.i_clk(tick), .i_in(), .o_out(w950107));
	wire w990107;
	torch #(1'b0) c990107 (.i_clk(tick), .i_in(), .o_out(w990107));
	wire w1030107;
	torch #(1'b0) c1030107 (.i_clk(tick), .i_in(), .o_out(w1030107));
	wire w1070107;
	torch #(1'b0) c1070107 (.i_clk(tick), .i_in(), .o_out(w1070107));
	wire w1110107;
	torch #(1'b0) c1110107 (.i_clk(tick), .i_in(), .o_out(w1110107));
	wire w1150107;
	torch #(1'b0) c1150107 (.i_clk(tick), .i_in(), .o_out(w1150107));
	wire w900109;
	torch #(1'b0) c900109 (.i_clk(tick), .i_in(), .o_out(w900109));
	wire w940109;
	torch #(1'b0) c940109 (.i_clk(tick), .i_in(), .o_out(w940109));
	wire w980109;
	torch #(1'b0) c980109 (.i_clk(tick), .i_in(), .o_out(w980109));
	wire w1020109;
	torch #(1'b1) c1020109 (.i_clk(tick), .i_in(), .o_out(w1020109));
	wire w1060109;
	torch #(1'b0) c1060109 (.i_clk(tick), .i_in(), .o_out(w1060109));
	wire w1100109;
	torch #(1'b0) c1100109 (.i_clk(tick), .i_in(), .o_out(w1100109));
	wire w1140109;
	torch #(1'b0) c1140109 (.i_clk(tick), .i_in(), .o_out(w1140109));
	wire w960111;
	torch #(1'b1) c960111 (.i_clk(tick), .i_in(), .o_out(w960111));
	wire w1000111;
	torch #(1'b1) c1000111 (.i_clk(tick), .i_in(), .o_out(w1000111));
	wire w1040111;
	torch #(1'b1) c1040111 (.i_clk(tick), .i_in(), .o_out(w1040111));
	wire w1080111;
	torch #(1'b1) c1080111 (.i_clk(tick), .i_in(), .o_out(w1080111));
	wire w900114;

	wire w940114;

	wire w980114;

	wire w1020114;

	wire w1060114;

	wire w1100114;

	wire w1140114;

	wire w440118;

	wire w620118;

	wire w910123;
	torch #(1'b0) c910123 (.i_clk(tick), .i_in(), .o_out(w910123));
	wire w950123;
	torch #(1'b0) c950123 (.i_clk(tick), .i_in(), .o_out(w950123));
	wire w990123;
	torch #(1'b0) c990123 (.i_clk(tick), .i_in(), .o_out(w990123));
	wire w1030123;
	torch #(1'b0) c1030123 (.i_clk(tick), .i_in(), .o_out(w1030123));
	wire w1070123;
	torch #(1'b0) c1070123 (.i_clk(tick), .i_in(), .o_out(w1070123));
	wire w1110123;
	torch #(1'b0) c1110123 (.i_clk(tick), .i_in(), .o_out(w1110123));
	wire w1150123;
	torch #(1'b0) c1150123 (.i_clk(tick), .i_in(), .o_out(w1150123));
	wire w900125;
	torch #(1'b0) c900125 (.i_clk(tick), .i_in(), .o_out(w900125));
	wire w940125;
	torch #(1'b0) c940125 (.i_clk(tick), .i_in(), .o_out(w940125));
	wire w980125;
	torch #(1'b0) c980125 (.i_clk(tick), .i_in(), .o_out(w980125));
	wire w1020125;
	torch #(1'b1) c1020125 (.i_clk(tick), .i_in(), .o_out(w1020125));
	wire w1060125;
	torch #(1'b0) c1060125 (.i_clk(tick), .i_in(), .o_out(w1060125));
	wire w1100125;
	torch #(1'b0) c1100125 (.i_clk(tick), .i_in(), .o_out(w1100125));
	wire w1140125;
	torch #(1'b0) c1140125 (.i_clk(tick), .i_in(), .o_out(w1140125));
	wire w960127;
	torch #(1'b1) c960127 (.i_clk(tick), .i_in(), .o_out(w960127));
	wire w1000127;
	torch #(1'b1) c1000127 (.i_clk(tick), .i_in(), .o_out(w1000127));
	wire w1040127;
	torch #(1'b1) c1040127 (.i_clk(tick), .i_in(), .o_out(w1040127));
	wire w1080127;
	torch #(1'b1) c1080127 (.i_clk(tick), .i_in(), .o_out(w1080127));
	wire w900130;

	wire w940130;

	wire w980130;

	wire w1020130;

	wire w1060130;

	wire w1100130;

	wire w1140130;

	wire w910139;
	torch #(1'b0) c910139 (.i_clk(tick), .i_in(), .o_out(w910139));
	wire w950139;
	torch #(1'b0) c950139 (.i_clk(tick), .i_in(), .o_out(w950139));
	wire w990139;
	torch #(1'b0) c990139 (.i_clk(tick), .i_in(), .o_out(w990139));
	wire w1030139;
	torch #(1'b0) c1030139 (.i_clk(tick), .i_in(), .o_out(w1030139));
	wire w1070139;
	torch #(1'b0) c1070139 (.i_clk(tick), .i_in(), .o_out(w1070139));
	wire w1110139;
	torch #(1'b0) c1110139 (.i_clk(tick), .i_in(), .o_out(w1110139));
	wire w1150139;
	torch #(1'b0) c1150139 (.i_clk(tick), .i_in(), .o_out(w1150139));
	wire w900141;
	torch #(1'b0) c900141 (.i_clk(tick), .i_in(), .o_out(w900141));
	wire w940141;
	torch #(1'b0) c940141 (.i_clk(tick), .i_in(), .o_out(w940141));
	wire w980141;
	torch #(1'b0) c980141 (.i_clk(tick), .i_in(), .o_out(w980141));
	wire w1020141;
	torch #(1'b1) c1020141 (.i_clk(tick), .i_in(), .o_out(w1020141));
	wire w1060141;
	torch #(1'b0) c1060141 (.i_clk(tick), .i_in(), .o_out(w1060141));
	wire w1100141;
	torch #(1'b0) c1100141 (.i_clk(tick), .i_in(), .o_out(w1100141));
	wire w1140141;
	torch #(1'b0) c1140141 (.i_clk(tick), .i_in(), .o_out(w1140141));
	wire w880144;
	assign outputs[19] = ();
	wire w900144;
	assign outputs[20] = ();
	wire w920144;
	assign outputs[21] = ();
	wire w940144;
	assign outputs[22] = ();
	wire w960144;
	assign outputs[23] = ();
	wire w980144;
	assign outputs[24] = ();
	wire w1000144;
	assign outputs[25] = ();
	wire w1020144;
	assign outputs[26] = ();
	wire w1040144;
	assign outputs[27] = ();
	wire w1060144;
	assign outputs[28] = ();
	wire w1080144;
	assign outputs[29] = ();
	wire w1100144;
	assign outputs[30] = ();
	wire w1120144;
	assign outputs[31] = ();
	wire w1140144;
	assign outputs[32] = ();
	wire w880145;
	repeater #(1, 1'b0, 0, 0) c880145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w880145));
	wire w900145;
	repeater #(1, 1'b0, 0, 0) c900145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w900145));
	wire w920145;
	repeater #(1, 1'b0, 0, 0) c920145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w920145));
	wire w940145;
	repeater #(1, 1'b0, 0, 0) c940145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w940145));
	wire w960145;
	repeater #(1, 1'b0, 0, 0) c960145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w960145));
	wire w980145;
	repeater #(1, 1'b0, 0, 0) c980145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w980145));
	wire w1000145;
	repeater #(1, 1'b1, 0, 0) c1000145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1000145));
	wire w1020145;
	repeater #(1, 1'b1, 0, 0) c1020145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1020145));
	wire w1040145;
	repeater #(1, 1'b0, 0, 0) c1040145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1040145));
	wire w1060145;
	repeater #(1, 1'b0, 0, 0) c1060145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060145));
	wire w1080145;
	repeater #(1, 1'b0, 0, 0) c1080145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1080145));
	wire w1100145;
	repeater #(1, 1'b0, 0, 0) c1100145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1100145));
	wire w1120145;
	repeater #(1, 1'b0, 0, 0) c1120145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1120145));
	wire w1140145;
	repeater #(1, 1'b0, 0, 0) c1140145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1140145));
	wire w890152;
	repeater #(2, 1'b1, 0, 0) c890152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w890152));
	wire w930152;
	repeater #(2, 1'b1, 0, 0) c930152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w930152));
	wire w970152;
	repeater #(2, 1'b1, 0, 0) c970152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w970152));
	wire w1010152;
	repeater #(2, 1'b0, 0, 0) c1010152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010152));
	wire w1050152;
	repeater #(2, 1'b1, 0, 0) c1050152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1050152));
	wire w1090152;
	repeater #(2, 1'b1, 0, 0) c1090152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1090152));
	wire w1130152;
	repeater #(2, 1'b1, 0, 0) c1130152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1130152));
	wire w870157;
	repeater #(1, 1'b1, 0, 0) c870157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w870157));
	wire w910157;
	repeater #(1, 1'b1, 0, 0) c910157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w910157));
	wire w950157;
	repeater #(1, 1'b1, 0, 0) c950157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w950157));
	wire w990157;
	repeater #(1, 1'b0, 0, 0) c990157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990157));
	wire w1030157;
	repeater #(1, 1'b1, 0, 0) c1030157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030157));
	wire w1070157;
	repeater #(1, 1'b1, 0, 0) c1070157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070157));
	wire w1110157;
	repeater #(1, 1'b1, 0, 0) c1110157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110157));
	wire w890158;

	wire w930158;

	wire w970158;

	wire w1010158;

	wire w1050158;

	wire w1090158;

	wire w1130158;

	wire w880159;

	wire w920159;

	wire w960159;

	wire w1000159;

	wire w1040159;

	wire w1080159;

	wire w1120159;

	wire w890160;
	torch #(1'b1) c890160 (.i_clk(tick), .i_in(), .o_out(w890160));
	wire w930160;
	torch #(1'b1) c930160 (.i_clk(tick), .i_in(), .o_out(w930160));
	wire w970160;
	torch #(1'b1) c970160 (.i_clk(tick), .i_in(), .o_out(w970160));
	wire w1010160;
	torch #(1'b1) c1010160 (.i_clk(tick), .i_in(), .o_out(w1010160));
	wire w1050160;
	torch #(1'b1) c1050160 (.i_clk(tick), .i_in(), .o_out(w1050160));
	wire w1090160;
	torch #(1'b1) c1090160 (.i_clk(tick), .i_in(), .o_out(w1090160));
	wire w1130160;
	torch #(1'b1) c1130160 (.i_clk(tick), .i_in(), .o_out(w1130160));
	wire w870161;
	repeater #(1, 1'b1, 0, 0) c870161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w870161));
	wire w910161;
	repeater #(1, 1'b1, 0, 0) c910161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w910161));
	wire w950161;
	repeater #(1, 1'b1, 0, 0) c950161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w950161));
	wire w990161;
	repeater #(1, 1'b1, 0, 0) c990161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990161));
	wire w1030161;
	repeater #(1, 1'b1, 0, 0) c1030161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030161));
	wire w1070161;
	repeater #(1, 1'b1, 0, 0) c1070161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070161));
	wire w1110161;
	repeater #(1, 1'b1, 0, 0) c1110161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110161));
	wire w870162;
	torch #(1'b0) c870162 (.i_clk(tick), .i_in(), .o_out(w870162));
	wire w890162;
	torch #(1'b0) c890162 (.i_clk(tick), .i_in(), .o_out(w890162));
	wire w910162;
	torch #(1'b0) c910162 (.i_clk(tick), .i_in(), .o_out(w910162));
	wire w930162;
	torch #(1'b0) c930162 (.i_clk(tick), .i_in(), .o_out(w930162));
	wire w950162;
	torch #(1'b0) c950162 (.i_clk(tick), .i_in(), .o_out(w950162));
	wire w970162;
	torch #(1'b0) c970162 (.i_clk(tick), .i_in(), .o_out(w970162));
	wire w990162;
	torch #(1'b0) c990162 (.i_clk(tick), .i_in(), .o_out(w990162));
	wire w1010162;
	torch #(1'b0) c1010162 (.i_clk(tick), .i_in(), .o_out(w1010162));
	wire w1030162;
	torch #(1'b0) c1030162 (.i_clk(tick), .i_in(), .o_out(w1030162));
	wire w1050162;
	torch #(1'b0) c1050162 (.i_clk(tick), .i_in(), .o_out(w1050162));
	wire w1070162;
	torch #(1'b0) c1070162 (.i_clk(tick), .i_in(), .o_out(w1070162));
	wire w1090162;
	torch #(1'b0) c1090162 (.i_clk(tick), .i_in(), .o_out(w1090162));
	wire w1110162;
	torch #(1'b0) c1110162 (.i_clk(tick), .i_in(), .o_out(w1110162));
	wire w1130162;
	torch #(1'b0) c1130162 (.i_clk(tick), .i_in(), .o_out(w1130162));
	wire w870164;

	wire w890164;
	repeater #(2, 1'b0, 0, 0) c890164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w890164));
	wire w910164;

	wire w930164;
	repeater #(2, 1'b0, 0, 0) c930164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w930164));
	wire w950164;

	wire w970164;
	repeater #(2, 1'b0, 0, 0) c970164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w970164));
	wire w990164;

	wire w1010164;
	repeater #(2, 1'b0, 0, 0) c1010164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010164));
	wire w1030164;

	wire w1050164;
	repeater #(2, 1'b0, 0, 0) c1050164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1050164));
	wire w1070164;

	wire w1090164;
	repeater #(2, 1'b0, 0, 0) c1090164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1090164));
	wire w1110164;

	wire w1130164;
	repeater #(2, 1'b0, 0, 0) c1130164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1130164));
	wire w1180165;
	repeater #(1, 1'b0, 0, 0) c1180165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1180165));
	wire w114140;

	wire w112142;

	wire w110144;

	wire w108146;

	wire w106148;

	wire w172152;
	repeater #(2, 1'b0, 0, 0) c172152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172152));
	wire w206152;
	repeater #(2, 1'b0, 0, 0) c206152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206152));
	wire w89154;
	torch #(1'b1) c89154 (.i_clk(tick), .i_in(), .o_out(w89154));
	wire w93154;
	torch #(1'b1) c93154 (.i_clk(tick), .i_in(), .o_out(w93154));
	wire w97154;
	torch #(1'b1) c97154 (.i_clk(tick), .i_in(), .o_out(w97154));
	wire w101154;
	torch #(1'b1) c101154 (.i_clk(tick), .i_in(), .o_out(w101154));
	wire w105154;
	torch #(1'b1) c105154 (.i_clk(tick), .i_in(), .o_out(w105154));
	wire w109154;
	torch #(1'b1) c109154 (.i_clk(tick), .i_in(), .o_out(w109154));
	wire w113154;
	torch #(1'b1) c113154 (.i_clk(tick), .i_in(), .o_out(w113154));
	wire w164154;
	torch #(1'b1) c164154 (.i_clk(tick), .i_in(), .o_out(w164154));
	wire w174154;
	repeater #(1, 1'b0, 0, 0) c174154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174154));
	wire w180154;
	torch #(1'b1) c180154 (.i_clk(tick), .i_in(), .o_out(w180154));
	wire w198154;
	torch #(1'b1) c198154 (.i_clk(tick), .i_in(), .o_out(w198154));
	wire w0155;
	repeater #(1, 1'b1, 0, 0) c0155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0155));
	wire w6155;
	torch #(1'b1) c6155 (.i_clk(tick), .i_in(), .o_out(w6155));
	wire w90157;
	repeater #(2, 1'b0, 0, 0) c90157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90157));
	wire w94157;
	repeater #(2, 1'b0, 0, 0) c94157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94157));
	wire w98157;
	repeater #(2, 1'b0, 0, 0) c98157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98157));
	wire w102157;
	repeater #(2, 1'b0, 0, 0) c102157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102157));
	wire w106157;
	repeater #(1, 1'b0, 0, 0) c106157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106157));
	wire w110157;
	repeater #(1, 1'b0, 0, 0) c110157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110157));
	wire w114157;
	repeater #(1, 1'b0, 0, 0) c114157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114157));
	wire w165157;
	repeater #(1, 1'b1, 0, 0) c165157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165157));
	wire w181157;
	repeater #(1, 1'b1, 0, 0) c181157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181157));
	wire w199157;
	repeater #(1, 1'b1, 0, 0) c199157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199157));
	wire w7158;
	repeater #(1, 1'b1, 0, 0) c7158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7158));
	wire w103158;
	repeater #(1, 1'b0, 0, 0) c103158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103158));
	wire w115158;
	repeater #(2, 1'b0, 0, 0) c115158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115158));
	wire w174158;
	repeater #(1, 1'b0, 0, 0) c174158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174158));
	wire w187158;

	wire w0159;
	repeater #(1, 1'b1, 0, 0) c0159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0159));
	wire w13159;

	wire w163159;

	wire w179159;

	wire w197159;

	wire w5160;

	wire w171160;

	wire w187160;

	wire w205160;

	wire w13161;

	wire w168161;

	wire w173161;

	wire w174161;

	wire w184161;

	wire w202161;

	wire w207161;

	wire w0162;

	wire w10162;

	wire w92163;
	repeater #(1, 1'b0, 0, 0) c92163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92163));
	wire w112163;
	repeater #(1, 1'b0, 0, 0) c112163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112163));
	wire w166163;

	wire w182163;

	wire w200163;

	wire w8164;

	wire w172164;

	wire w173164;

	wire w206164;

	wire w207164;

	wire w158165;

	wire w192165;

	wire w29166;
	repeater #(1, 1'b1, 0, 0) c29166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29166));
	wire w31166;
	repeater #(2, 1'b0, 0, 0) c31166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31166));
	wire w33166;
	repeater #(2, 1'b0, 0, 0) c33166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33166));
	wire w37166;
	repeater #(2, 1'b1, 0, 0) c37166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37166));
	wire w39166;
	repeater #(2, 1'b0, 0, 0) c39166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39166));
	wire w41166;
	repeater #(1, 1'b1, 0, 0) c41166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41166));
	wire w61166;
	repeater #(1, 1'b1, 0, 0) c61166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61166));
	wire w63166;
	repeater #(2, 1'b1, 0, 0) c63166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63166));
	wire w65166;
	repeater #(2, 1'b0, 0, 0) c65166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65166));
	wire w69166;
	repeater #(2, 1'b1, 0, 0) c69166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69166));
	wire w71166;
	repeater #(2, 1'b1, 0, 0) c71166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71166));
	wire w73166;
	repeater #(1, 1'b1, 0, 0) c73166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73166));
	wire w26167;
	repeater #(1, 1'b1, 0, 0) c26167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26167));
	wire w76167;
	repeater #(1, 1'b1, 0, 0) c76167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76167));
	wire w159167;
	repeater #(1, 1'b1, 0, 0) c159167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159167));
	wire w163167;
	repeater #(1, 1'b1, 0, 0) c163167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163167));
	wire w167167;
	repeater #(1, 1'b1, 0, 0) c167167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167167));
	wire w171167;
	repeater #(1, 1'b0, 0, 0) c171167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171167));
	wire w175167;
	repeater #(1, 1'b1, 0, 0) c175167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175167));
	wire w179167;
	repeater #(1, 1'b1, 0, 0) c179167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179167));
	wire w183167;
	repeater #(1, 1'b1, 0, 0) c183167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183167));
	wire w193167;
	repeater #(1, 1'b1, 0, 0) c193167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193167));
	wire w197167;
	repeater #(1, 1'b1, 0, 0) c197167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197167));
	wire w201167;
	repeater #(1, 1'b1, 0, 0) c201167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201167));
	wire w205167;
	repeater #(1, 1'b1, 0, 0) c205167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205167));
	wire w1168;
	repeater #(1, 1'b1, 0, 0) c1168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1168));
	wire w5168;
	repeater #(1, 1'b1, 0, 0) c5168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5168));
	wire w9168;
	repeater #(1, 1'b1, 0, 0) c9168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9168));
	wire w36168;

	wire w66168;

	wire w28169;

	wire w32169;

	wire w35169;

	wire w37169;

	wire w40169;

	wire w62169;

	wire w65169;

	wire w67169;

	wire w70169;

	wire w74169;

	wire w27170;

	wire w29170;

	wire w31170;

	wire w33170;

	wire w36170;

	wire w39170;

	wire w41170;

	wire w61170;

	wire w63170;

	wire w66170;

	wire w69170;

	wire w71170;

	wire w73170;

	wire w75170;

	wire w32171;

	wire w70171;

	wire w28172;

	wire w32172;

	wire w33172;

	wire w37172;

	wire w39172;

	wire w41172;

	wire w61172;

	wire w63172;

	wire w65172;

	wire w69172;

	wire w70172;

	wire w74172;

	wire w27174;

	wire w33174;

	wire w69174;

	wire w75174;

	wire w23175;
	repeater #(1, 1'b1, 0, 0) c23175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23175));
	wire w28175;
	repeater #(1, 1'b1, 0, 0) c28175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28175));
	wire w33175;
	repeater #(1, 1'b1, 0, 0) c33175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33175));
	wire w69175;
	repeater #(1, 1'b0, 0, 0) c69175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69175));
	wire w74175;
	repeater #(1, 1'b1, 0, 0) c74175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74175));
	wire w79175;
	repeater #(1, 1'b1, 0, 0) c79175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79175));
	wire w166176;

	wire w200176;

	wire w164177;
	repeater #(1, 1'b1, 0, 0) c164177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164177));
	wire w198177;
	repeater #(1, 1'b1, 0, 0) c198177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198177));
	wire w155178;
	repeater #(1, 1'b1, 0, 0) c155178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155178));
	wire w171178;
	repeater #(1, 1'b1, 0, 0) c171178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171178));
	wire w189178;
	repeater #(1, 1'b1, 0, 0) c189178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189178));
	wire w205178;
	repeater #(1, 1'b1, 0, 0) c205178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205178));
	wire w22179;

	wire w23179;
	repeater #(1, 1'b0, 0, 0) c23179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23179));
	wire w27179;

	wire w28179;
	repeater #(1, 1'b0, 0, 0) c28179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28179));
	wire w32179;

	wire w33179;
	repeater #(1, 1'b0, 0, 0) c33179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33179));
	wire w69179;
	repeater #(1, 1'b0, 0, 0) c69179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69179));
	wire w70179;

	wire w74179;
	repeater #(1, 1'b1, 0, 0) c74179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74179));
	wire w75179;

	wire w79179;
	repeater #(1, 1'b1, 0, 0) c79179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79179));
	wire w80179;

	wire w92179;
	repeater #(1, 1'b0, 0, 0) c92179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92179));
	wire w112179;
	repeater #(1, 1'b0, 0, 0) c112179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112179));
	wire w166179;

	wire w182179;

	wire w200179;

	wire w8180;

	wire w158180;

	wire w174180;

	wire w192180;

	wire w0181;

	wire w155181;

	wire w156181;

	wire w161181;

	wire w169181;

	wire w171181;

	wire w172181;

	wire w177181;

	wire w185181;

	wire w189181;

	wire w190181;

	wire w195181;

	wire w203181;

	wire w205181;

	wire w206181;

	wire w3182;

	wire w11182;

	wire w182182;

	wire w8183;

	wire w23183;
	repeater #(2, 1'b0, 0, 0) c23183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23183));
	wire w28183;
	repeater #(2, 1'b0, 0, 0) c28183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28183));
	wire w33183;
	repeater #(2, 1'b0, 0, 0) c33183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33183));
	wire w69183;
	repeater #(2, 1'b0, 0, 0) c69183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69183));
	wire w74183;
	repeater #(2, 1'b1, 0, 0) c74183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74183));
	wire w79183;
	repeater #(2, 1'b1, 0, 0) c79183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79183));
	wire w163183;

	wire w164183;

	wire w179183;

	wire w180183;

	wire w197183;

	wire w198183;

	wire w5184;

	wire w6184;

	wire w155185;

	wire w156185;

	wire w169185;

	wire w171185;

	wire w172185;

	wire w185185;

	wire w189185;

	wire w190185;

	wire w203185;

	wire w205185;

	wire w206185;

	wire w11186;

	wire w49186;

	wire w40187;
	repeater #(1, 1'b0, 0, 0) c40187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40187));
	wire w62187;
	repeater #(1, 1'b0, 0, 0) c62187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62187));
	wire w166187;
	torch #(1'b1) c166187 (.i_clk(tick), .i_in(), .o_out(w166187));
	wire w167187;

	wire w182187;
	torch #(1'b1) c182187 (.i_clk(tick), .i_in(), .o_out(w182187));
	wire w183187;

	wire w200187;
	torch #(1'b1) c200187 (.i_clk(tick), .i_in(), .o_out(w200187));
	wire w201187;

	wire w8188;
	torch #(1'b1) c8188 (.i_clk(tick), .i_in(), .o_out(w8188));
	wire w9188;

	wire w51188;

	wire w167188;

	wire w169188;

	wire w183188;

	wire w185188;

	wire w201188;

	wire w203188;

	wire w9189;

	wire w11189;

	wire w22189;

	wire w23189;

	wire w52189;

	wire w79189;

	wire w80189;

	wire w26190;
	repeater #(2, 1'b0, 0, 0) c26190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26190));
	wire w27190;
	repeater #(2, 1'b0, 0, 0) c27190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27190));
	wire w29190;

	wire w43190;
	repeater #(1, 1'b0, 0, 0) c43190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43190));
	wire w44190;

	wire w52190;
	repeater #(1, 1'b1, 0, 0) c52190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52190));
	wire w58190;

	wire w59190;
	repeater #(1, 1'b1, 0, 0) c59190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59190));
	wire w73190;

	wire w75190;
	repeater #(2, 1'b0, 0, 0) c75190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75190));
	wire w76190;
	repeater #(2, 1'b0, 0, 0) c76190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76190));
	wire w169190;

	wire w170190;

	wire w171190;

	wire w185190;

	wire w186190;

	wire w187190;

	wire w203190;

	wire w204190;

	wire w205190;

	wire w11191;

	wire w12191;

	wire w13191;

	wire w27191;

	wire w29191;
	repeater #(1, 1'b1, 0, 0) c29191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29191));
	wire w40191;

	wire w41191;

	wire w61191;

	wire w62191;

	wire w73191;
	repeater #(1, 1'b1, 0, 0) c73191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73191));
	wire w75191;

	wire w164191;

	wire w165191;

	wire w171191;

	wire w180191;

	wire w181191;

	wire w187191;

	wire w198191;

	wire w199191;

	wire w205191;

	wire w6192;

	wire w7192;

	wire w13192;

	wire w23192;

	wire w27192;

	wire w51192;

	wire w52192;

	wire w75192;

	wire w79192;

	wire w23193;

	wire w25193;
	repeater #(1, 1'b0, 0, 0) c25193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25193));
	wire w30193;

	wire w34193;

	wire w40193;
	repeater #(1, 1'b0, 0, 0) c40193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40193));
	wire w48193;

	wire w49193;
	repeater #(1, 1'b1, 0, 0) c49193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49193));
	wire w62193;
	repeater #(1, 1'b0, 0, 0) c62193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62193));
	wire w68193;

	wire w72193;

	wire w77193;
	repeater #(1, 1'b0, 0, 0) c77193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77193));
	wire w79193;

	wire w161193;
	torch #(1'b0) c161193 (.i_clk(tick), .i_in(), .o_out(w161193));
	wire w169193;
	repeater #(1, 1'b0, 0, 0) c169193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169193));
	wire w171193;
	torch #(1'b0) c171193 (.i_clk(tick), .i_in(), .o_out(w171193));
	wire w177193;
	torch #(1'b0) c177193 (.i_clk(tick), .i_in(), .o_out(w177193));
	wire w185193;
	repeater #(1, 1'b0, 0, 0) c185193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185193));
	wire w187193;
	torch #(1'b0) c187193 (.i_clk(tick), .i_in(), .o_out(w187193));
	wire w195193;
	torch #(1'b0) c195193 (.i_clk(tick), .i_in(), .o_out(w195193));
	wire w203193;
	repeater #(1, 1'b0, 0, 0) c203193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203193));
	wire w205193;
	torch #(1'b0) c205193 (.i_clk(tick), .i_in(), .o_out(w205193));
	wire w3194;
	torch #(1'b0) c3194 (.i_clk(tick), .i_in(), .o_out(w3194));
	wire w11194;
	repeater #(1, 1'b0, 0, 0) c11194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11194));
	wire w13194;
	torch #(1'b0) c13194 (.i_clk(tick), .i_in(), .o_out(w13194));
	wire w30194;

	wire w32194;
	repeater #(1, 1'b1, 0, 0) c32194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32194));
	wire w33194;

	wire w40194;

	wire w57194;

	wire w62194;

	wire w69194;

	wire w70194;
	repeater #(1, 1'b1, 0, 0) c70194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70194));
	wire w72194;

	wire w26195;

	wire w41195;

	wire w45195;
	repeater #(1, 1'b0, 0, 0) c45195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45195));
	wire w58195;
	repeater #(2, 1'b0, 0, 0) c58195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58195));
	wire w61195;

	wire w76195;

	wire w92195;
	repeater #(1, 1'b0, 0, 0) c92195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92195));
	wire w112195;
	repeater #(1, 1'b0, 0, 0) c112195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112195));
	wire w173195;
	repeater #(1, 1'b1, 0, 0) c173195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173195));
	wire w207195;
	repeater #(1, 1'b1, 0, 0) c207195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207195));
	wire w23196;

	wire w24196;
	repeater #(1, 1'b1, 0, 0) c24196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24196));
	wire w31196;
	repeater #(2, 1'b1, 0, 0) c31196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31196));
	wire w44196;
	assign outputs[33] = ();
	wire w71196;
	repeater #(2, 1'b1, 0, 0) c71196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71196));
	wire w78196;
	repeater #(1, 1'b0, 0, 0) c78196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78196));
	wire w79196;

	wire w170197;
	torch #(1'b1) c170197 (.i_clk(tick), .i_in(), .o_out(w170197));
	wire w186197;
	torch #(1'b1) c186197 (.i_clk(tick), .i_in(), .o_out(w186197));
	wire w204197;
	torch #(1'b1) c204197 (.i_clk(tick), .i_in(), .o_out(w204197));
	wire w12198;
	torch #(1'b1) c12198 (.i_clk(tick), .i_in(), .o_out(w12198));
	wire w162199;
	torch #(1'b1) c162199 (.i_clk(tick), .i_in(), .o_out(w162199));
	wire w178199;
	torch #(1'b1) c178199 (.i_clk(tick), .i_in(), .o_out(w178199));
	wire w196199;
	torch #(1'b1) c196199 (.i_clk(tick), .i_in(), .o_out(w196199));
	wire w41100;
	torch #(1'b1) c41100 (.i_clk(tick), .i_in(), .o_out(w41100));
	wire w1691100;
	repeater #(1, 1'b0, 0, 0) c1691100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1691100));
	wire w1851100;
	repeater #(1, 1'b0, 0, 0) c1851100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1851100));
	wire w2031100;
	repeater #(1, 1'b0, 0, 0) c2031100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2031100));
	wire w111101;
	repeater #(1, 1'b0, 0, 0) c111101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111101));
	wire w1631101;
	repeater #(1, 1'b0, 0, 0) c1631101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1631101));
	wire w1791101;
	repeater #(1, 1'b0, 0, 0) c1791101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1791101));
	wire w1971101;
	repeater #(1, 1'b0, 0, 0) c1971101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1971101));
	wire w51102;
	repeater #(1, 1'b0, 0, 0) c51102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51102));
	wire w921111;
	repeater #(1, 1'b0, 0, 0) c921111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w921111));
	wire w1121111;
	repeater #(1, 1'b0, 0, 0) c1121111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121111));
	wire w501118;

	wire w511118;
	repeater #(1, 1'b0, 0, 0) c511118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w511118));
	wire w521119;
	repeater #(1, 1'b0, 0, 0) c521119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w521119));
	wire w551119;
	repeater #(2, 1'b0, 0, 0) c551119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w551119));
	wire w471120;
	repeater #(1, 1'b0, 0, 0) c471120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w471120));
	wire w601120;
	repeater #(2, 1'b0, 0, 0) c601120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w601120));
	wire w461121;
	assign outputs[34] = ();
	wire w491121;

	wire w581121;

	wire w491122;

	wire w581122;

	wire w471123;
	repeater #(1, 1'b0, 0, 0) c471123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w471123));
	wire w601123;
	repeater #(1, 1'b0, 0, 0) c601123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w601123));
	wire w921127;
	repeater #(1, 1'b0, 0, 0) c921127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w921127));
	wire w1121127;
	repeater #(1, 1'b0, 0, 0) c1121127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121127));
	wire w73012;
	torch #(1'b1) c73012 (.i_clk(tick), .i_in(), .o_out(w73012));
	wire w77012;
	torch #(1'b1) c77012 (.i_clk(tick), .i_in(), .o_out(w77012));
	wire w81012;
	torch #(1'b1) c81012 (.i_clk(tick), .i_in(), .o_out(w81012));
	wire w85012;
	torch #(1'b0) c85012 (.i_clk(tick), .i_in(), .o_out(w85012));
	wire w89012;
	torch #(1'b1) c89012 (.i_clk(tick), .i_in(), .o_out(w89012));
	wire w93012;
	torch #(1'b1) c93012 (.i_clk(tick), .i_in(), .o_out(w93012));
	wire w97012;
	torch #(1'b1) c97012 (.i_clk(tick), .i_in(), .o_out(w97012));
	wire w73016;
	torch #(1'b1) c73016 (.i_clk(tick), .i_in(), .o_out(w73016));
	wire w77016;
	torch #(1'b1) c77016 (.i_clk(tick), .i_in(), .o_out(w77016));
	wire w81016;
	torch #(1'b1) c81016 (.i_clk(tick), .i_in(), .o_out(w81016));
	wire w85016;
	torch #(1'b1) c85016 (.i_clk(tick), .i_in(), .o_out(w85016));
	wire w89016;
	torch #(1'b1) c89016 (.i_clk(tick), .i_in(), .o_out(w89016));
	wire w93016;
	torch #(1'b1) c93016 (.i_clk(tick), .i_in(), .o_out(w93016));
	wire w97016;
	torch #(1'b1) c97016 (.i_clk(tick), .i_in(), .o_out(w97016));
	wire w72024;
	torch #(1'b1) c72024 (.i_clk(tick), .i_in(), .o_out(w72024));
	wire w76024;
	torch #(1'b1) c76024 (.i_clk(tick), .i_in(), .o_out(w76024));
	wire w80024;
	torch #(1'b1) c80024 (.i_clk(tick), .i_in(), .o_out(w80024));
	wire w84024;
	torch #(1'b1) c84024 (.i_clk(tick), .i_in(), .o_out(w84024));
	wire w88024;
	torch #(1'b1) c88024 (.i_clk(tick), .i_in(), .o_out(w88024));
	wire w92024;
	torch #(1'b1) c92024 (.i_clk(tick), .i_in(), .o_out(w92024));
	wire w96024;
	torch #(1'b1) c96024 (.i_clk(tick), .i_in(), .o_out(w96024));
	wire w73057;
	repeater #(1, 1'b0, 0, 0) c73057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73057));
	wire w77057;
	repeater #(1, 1'b0, 0, 0) c77057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77057));
	wire w81057;
	repeater #(1, 1'b0, 0, 0) c81057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81057));
	wire w85057;
	repeater #(1, 1'b0, 0, 0) c85057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85057));
	wire w89057;
	repeater #(1, 1'b0, 0, 0) c89057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89057));
	wire w93057;
	repeater #(1, 1'b0, 0, 0) c93057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93057));
	wire w97057;
	repeater #(1, 1'b0, 0, 0) c97057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97057));
	wire w73060;
	torch #(1'b1) c73060 (.i_clk(tick), .i_in(), .o_out(w73060));
	wire w77060;
	torch #(1'b1) c77060 (.i_clk(tick), .i_in(), .o_out(w77060));
	wire w81060;
	torch #(1'b1) c81060 (.i_clk(tick), .i_in(), .o_out(w81060));
	wire w85060;
	torch #(1'b1) c85060 (.i_clk(tick), .i_in(), .o_out(w85060));
	wire w89060;
	torch #(1'b1) c89060 (.i_clk(tick), .i_in(), .o_out(w89060));
	wire w93060;
	torch #(1'b1) c93060 (.i_clk(tick), .i_in(), .o_out(w93060));
	wire w97060;
	torch #(1'b1) c97060 (.i_clk(tick), .i_in(), .o_out(w97060));
	wire w84063;
	repeater #(1, 1'b0, 0, 0) c84063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84063));
	wire w86063;
	repeater #(1, 1'b1, 0, 0) c86063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86063));
	wire w88063;
	repeater #(1, 1'b1, 0, 0) c88063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88063));
	wire w90063;
	repeater #(1, 1'b1, 0, 0) c90063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90063));
	wire w92063;
	repeater #(1, 1'b1, 0, 0) c92063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92063));
	wire w94063;
	repeater #(1, 1'b1, 0, 0) c94063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94063));
	wire w96063;
	repeater #(1, 1'b1, 0, 0) c96063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96063));
	wire w98063;
	repeater #(1, 1'b1, 0, 0) c98063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98063));
	wire w82065;
	repeater #(1, 1'b1, 0, 0) c82065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82065));
	wire w80067;
	repeater #(1, 1'b1, 0, 0) c80067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80067));
	wire w78069;
	repeater #(1, 1'b1, 0, 0) c78069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78069));
	wire w76071;
	repeater #(1, 1'b1, 0, 0) c76071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76071));
	wire w74073;
	repeater #(1, 1'b1, 0, 0) c74073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74073));
	wire w72075;
	repeater #(1, 1'b1, 0, 0) c72075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72075));
	wire w170080;
	torch #(1'b1) c170080 (.i_clk(tick), .i_in(), .o_out(w170080));
	wire w204080;
	repeater #(1, 1'b1, 0, 0) c204080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204080));
	wire w30081;
	torch #(1'b1) c30081 (.i_clk(tick), .i_in(), .o_out(w30081));
	wire w64081;
	repeater #(1, 1'b1, 0, 0) c64081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64081));
	wire w168082;
	repeater #(1, 1'b1, 0, 0) c168082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168082));
	wire w202082;
	repeater #(1, 1'b1, 0, 0) c202082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202082));
	wire w28083;
	repeater #(1, 1'b1, 0, 0) c28083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28083));
	wire w62083;
	repeater #(1, 1'b1, 0, 0) c62083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62083));
	wire w98084;
	repeater #(1, 1'b1, 0, 0) c98084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98084));
	wire w166084;
	torch #(1'b1) c166084 (.i_clk(tick), .i_in(), .o_out(w166084));
	wire w200084;
	repeater #(1, 1'b1, 0, 0) c200084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200084));
	wire w26085;
	torch #(1'b1) c26085 (.i_clk(tick), .i_in(), .o_out(w26085));
	wire w60085;
	repeater #(1, 1'b1, 0, 0) c60085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60085));
	wire w96086;
	repeater #(1, 1'b1, 0, 0) c96086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96086));
	wire w164086;
	repeater #(1, 1'b1, 0, 0) c164086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164086));
	wire w198086;
	repeater #(1, 1'b1, 0, 0) c198086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198086));
	wire w24087;
	repeater #(1, 1'b1, 0, 0) c24087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24087));
	wire w58087;
	repeater #(1, 1'b1, 0, 0) c58087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58087));
	wire w94088;
	repeater #(1, 1'b1, 0, 0) c94088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94088));
	wire w162088;
	torch #(1'b1) c162088 (.i_clk(tick), .i_in(), .o_out(w162088));
	wire w196088;
	repeater #(1, 1'b1, 0, 0) c196088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196088));
	wire w22089;
	torch #(1'b1) c22089 (.i_clk(tick), .i_in(), .o_out(w22089));
	wire w56089;
	repeater #(1, 1'b1, 0, 0) c56089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56089));
	wire w92090;
	repeater #(1, 1'b1, 0, 0) c92090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92090));
	wire w160090;
	repeater #(1, 1'b1, 0, 0) c160090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160090));
	wire w194090;
	repeater #(1, 1'b1, 0, 0) c194090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194090));
	wire w20091;
	repeater #(1, 1'b1, 0, 0) c20091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20091));
	wire w54091;
	repeater #(1, 1'b1, 0, 0) c54091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54091));
	wire w144091;
	repeater #(1, 1'b1, 0, 0) c144091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144091));
	wire w146091;
	torch #(1'b1) c146091 (.i_clk(tick), .i_in(), .o_out(w146091));
	wire w148091;
	repeater #(1, 1'b1, 0, 0) c148091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148091));
	wire w150091;
	torch #(1'b1) c150091 (.i_clk(tick), .i_in(), .o_out(w150091));
	wire w152091;
	repeater #(1, 1'b1, 0, 0) c152091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152091));
	wire w154091;
	torch #(1'b1) c154091 (.i_clk(tick), .i_in(), .o_out(w154091));
	wire w156091;
	repeater #(1, 1'b0, 0, 0) c156091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156091));
	wire w158091;
	torch #(1'b1) c158091 (.i_clk(tick), .i_in(), .o_out(w158091));
	wire w178091;
	repeater #(1, 1'b1, 0, 0) c178091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178091));
	wire w180091;
	repeater #(1, 1'b1, 0, 0) c180091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180091));
	wire w182091;
	repeater #(1, 1'b1, 0, 0) c182091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182091));
	wire w184091;
	repeater #(1, 1'b1, 0, 0) c184091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184091));
	wire w186091;
	repeater #(1, 1'b1, 0, 0) c186091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186091));
	wire w188091;
	repeater #(1, 1'b1, 0, 0) c188091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188091));
	wire w190091;
	repeater #(1, 1'b0, 0, 0) c190091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190091));
	wire w192091;
	repeater #(1, 1'b1, 0, 0) c192091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192091));
	wire w6092;
	torch #(1'b1) c6092 (.i_clk(tick), .i_in(), .o_out(w6092));
	wire w10092;
	torch #(1'b1) c10092 (.i_clk(tick), .i_in(), .o_out(w10092));
	wire w14092;
	torch #(1'b1) c14092 (.i_clk(tick), .i_in(), .o_out(w14092));
	wire w18092;
	torch #(1'b1) c18092 (.i_clk(tick), .i_in(), .o_out(w18092));
	wire w38092;
	repeater #(1, 1'b1, 0, 0) c38092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38092));
	wire w40092;
	repeater #(1, 1'b1, 0, 0) c40092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40092));
	wire w42092;
	repeater #(1, 1'b1, 0, 0) c42092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42092));
	wire w44092;
	repeater #(1, 1'b1, 0, 0) c44092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44092));
	wire w46092;
	repeater #(1, 1'b1, 0, 0) c46092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46092));
	wire w48092;
	repeater #(1, 1'b1, 0, 0) c48092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48092));
	wire w50092;
	repeater #(1, 1'b0, 0, 0) c50092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50092));
	wire w52092;
	repeater #(1, 1'b1, 0, 0) c52092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52092));
	wire w90092;
	repeater #(1, 1'b1, 0, 0) c90092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90092));
	wire w5093;
	repeater #(1, 1'b1, 0, 0) c5093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5093));
	wire w9093;
	repeater #(1, 1'b1, 0, 0) c9093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9093));
	wire w13093;
	repeater #(1, 1'b1, 0, 0) c13093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13093));
	wire w17093;
	repeater #(1, 1'b0, 0, 0) c17093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17093));
	wire w76093;
	repeater #(1, 1'b1, 0, 0) c76093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76093));
	wire w78093;
	repeater #(1, 1'b1, 0, 0) c78093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78093));
	wire w80093;
	repeater #(1, 1'b1, 0, 0) c80093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80093));
	wire w82093;
	repeater #(1, 1'b1, 0, 0) c82093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82093));
	wire w84093;
	repeater #(1, 1'b0, 0, 0) c84093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84093));
	wire w86093;
	repeater #(1, 1'b1, 0, 0) c86093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86093));
	wire w88093;
	repeater #(1, 1'b1, 0, 0) c88093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88093));
	wire w6095;
	torch #(1'b1) c6095 (.i_clk(tick), .i_in(), .o_out(w6095));
	wire w10095;
	torch #(1'b1) c10095 (.i_clk(tick), .i_in(), .o_out(w10095));
	wire w14095;
	torch #(1'b1) c14095 (.i_clk(tick), .i_in(), .o_out(w14095));
	wire w18095;
	torch #(1'b0) c18095 (.i_clk(tick), .i_in(), .o_out(w18095));
	wire w22095;
	torch #(1'b1) c22095 (.i_clk(tick), .i_in(), .o_out(w22095));
	wire w26095;
	torch #(1'b1) c26095 (.i_clk(tick), .i_in(), .o_out(w26095));
	wire w30095;
	torch #(1'b1) c30095 (.i_clk(tick), .i_in(), .o_out(w30095));
	wire w40095;
	torch #(1'b1) c40095 (.i_clk(tick), .i_in(), .o_out(w40095));
	wire w44095;
	torch #(1'b1) c44095 (.i_clk(tick), .i_in(), .o_out(w44095));
	wire w48095;
	torch #(1'b1) c48095 (.i_clk(tick), .i_in(), .o_out(w48095));
	wire w52095;
	torch #(1'b1) c52095 (.i_clk(tick), .i_in(), .o_out(w52095));
	wire w56095;
	torch #(1'b1) c56095 (.i_clk(tick), .i_in(), .o_out(w56095));
	wire w60095;
	torch #(1'b1) c60095 (.i_clk(tick), .i_in(), .o_out(w60095));
	wire w64095;
	torch #(1'b1) c64095 (.i_clk(tick), .i_in(), .o_out(w64095));
	wire w144095;
	repeater #(2, 1'b1, 0, 0) c144095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144095));
	wire w148095;
	repeater #(2, 1'b1, 0, 0) c148095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148095));
	wire w152095;
	repeater #(2, 1'b1, 0, 0) c152095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152095));
	wire w168095;
	repeater #(2, 1'b1, 0, 0) c168095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168095));
	wire w178095;
	repeater #(2, 1'b1, 0, 0) c178095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178095));
	wire w182095;
	repeater #(2, 1'b1, 0, 0) c182095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182095));
	wire w186095;
	repeater #(2, 1'b1, 0, 0) c186095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186095));
	wire w202095;
	repeater #(2, 1'b1, 0, 0) c202095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202095));
	wire w11097;
	torch #(1'b1) c11097 (.i_clk(tick), .i_in(), .o_out(w11097));
	wire w15097;
	torch #(1'b1) c15097 (.i_clk(tick), .i_in(), .o_out(w15097));
	wire w19097;
	torch #(1'b1) c19097 (.i_clk(tick), .i_in(), .o_out(w19097));
	wire w23097;
	torch #(1'b1) c23097 (.i_clk(tick), .i_in(), .o_out(w23097));
	wire w47097;
	torch #(1'b0) c47097 (.i_clk(tick), .i_in(), .o_out(w47097));
	wire w51097;
	torch #(1'b0) c51097 (.i_clk(tick), .i_in(), .o_out(w51097));
	wire w55097;
	torch #(1'b0) c55097 (.i_clk(tick), .i_in(), .o_out(w55097));
	wire w59097;
	torch #(1'b0) c59097 (.i_clk(tick), .i_in(), .o_out(w59097));
	wire w144097;
	torch #(1'b1) c144097 (.i_clk(tick), .i_in(), .o_out(w144097));
	wire w154097;
	repeater #(1, 1'b1, 0, 0) c154097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154097));
	wire w160097;
	torch #(1'b1) c160097 (.i_clk(tick), .i_in(), .o_out(w160097));
	wire w170097;
	repeater #(1, 1'b1, 0, 0) c170097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170097));
	wire w178097;
	torch #(1'b1) c178097 (.i_clk(tick), .i_in(), .o_out(w178097));
	wire w188097;
	repeater #(1, 1'b1, 0, 0) c188097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188097));
	wire w194097;
	torch #(1'b1) c194097 (.i_clk(tick), .i_in(), .o_out(w194097));
	wire w204097;
	repeater #(1, 1'b1, 0, 0) c204097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204097));
	wire w1610100;
	repeater #(1, 1'b1, 0, 0) c1610100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610100));
	wire w1950100;
	repeater #(1, 1'b1, 0, 0) c1950100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950100));
	wire w1540101;
	repeater #(1, 1'b1, 0, 0) c1540101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540101));
	wire w1700101;
	repeater #(1, 1'b1, 0, 0) c1700101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1700101));
	wire w1880101;
	repeater #(1, 1'b1, 0, 0) c1880101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1880101));
	wire w2040101;
	repeater #(1, 1'b1, 0, 0) c2040101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040101));
	wire w1430102;

	wire w1590102;

	wire w1770102;

	wire w1930102;

	wire w740103;
	repeater #(1, 1'b1, 0, 0) c740103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w740103));
	wire w780103;
	repeater #(1, 1'b1, 0, 0) c780103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w780103));
	wire w820103;
	repeater #(1, 1'b1, 0, 0) c820103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w820103));
	wire w860103;
	repeater #(1, 1'b0, 0, 0) c860103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w860103));
	wire w900103;
	repeater #(1, 1'b1, 0, 0) c900103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w900103));
	wire w940103;
	repeater #(1, 1'b1, 0, 0) c940103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w940103));
	wire w980103;
	repeater #(1, 1'b1, 0, 0) c980103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w980103));
	wire w1510103;

	wire w1670103;

	wire w1850103;

	wire w2010103;

	wire w1480104;

	wire w1530104;

	wire w1540104;

	wire w1640104;

	wire w1690104;

	wire w1700104;

	wire w1820104;

	wire w1870104;

	wire w1880104;

	wire w1980104;

	wire w2030104;

	wire w2040104;

	wire w1430105;

	wire w1770105;

	wire w1460106;

	wire w1620106;

	wire w1800106;

	wire w1960106;

	wire w1010107;
	repeater #(1, 1'b0, 0, 0) c1010107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010107));
	wire w1520107;

	wire w1530107;

	wire w1680107;

	wire w1690107;

	wire w1860107;

	wire w1870107;

	wire w2020107;

	wire w2030107;

	wire w1620108;

	wire w1660108;

	wire w1960108;

	wire w2000108;

	wire w710109;
	repeater #(1, 1'b0, 0, 0) c710109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710109));
	wire w800112;
	torch #(1'b1) c800112 (.i_clk(tick), .i_in(), .o_out(w800112));
	wire w840112;
	torch #(1'b1) c840112 (.i_clk(tick), .i_in(), .o_out(w840112));
	wire w880112;
	torch #(1'b1) c880112 (.i_clk(tick), .i_in(), .o_out(w880112));
	wire w920112;
	torch #(1'b1) c920112 (.i_clk(tick), .i_in(), .o_out(w920112));
	wire w1430112;

	wire w1440112;

	wire w1470112;

	wire w1480112;

	wire w1510112;

	wire w1520112;

	wire w1550112;

	wire w1560112;

	wire w1590112;

	wire w1600112;

	wire w1630112;

	wire w1640112;

	wire w1670112;

	wire w1680112;

	wire w1770112;

	wire w1780112;

	wire w1810112;

	wire w1820112;

	wire w1850112;

	wire w1860112;

	wire w1890112;

	wire w1900112;

	wire w1930112;

	wire w1940112;

	wire w1970112;

	wire w1980112;

	wire w2010112;

	wire w2020112;

	wire w1440114;

	wire w1480114;

	wire w1520114;

	wire w1560114;

	wire w1600114;

	wire w1640114;

	wire w1680114;

	wire w1780114;

	wire w1820114;

	wire w1860114;

	wire w1900114;

	wire w1940114;

	wire w1980114;

	wire w2020114;

	wire w730116;
	torch #(1'b0) c730116 (.i_clk(tick), .i_in(), .o_out(w730116));
	wire w770116;
	torch #(1'b0) c770116 (.i_clk(tick), .i_in(), .o_out(w770116));
	wire w810116;
	torch #(1'b0) c810116 (.i_clk(tick), .i_in(), .o_out(w810116));
	wire w850116;
	torch #(1'b1) c850116 (.i_clk(tick), .i_in(), .o_out(w850116));
	wire w890116;
	torch #(1'b0) c890116 (.i_clk(tick), .i_in(), .o_out(w890116));
	wire w930116;
	torch #(1'b0) c930116 (.i_clk(tick), .i_in(), .o_out(w930116));
	wire w970116;
	torch #(1'b0) c970116 (.i_clk(tick), .i_in(), .o_out(w970116));
	wire w1420117;

	wire w1460117;

	wire w1500117;

	wire w1540117;

	wire w1760117;

	wire w1800117;

	wire w1840117;

	wire w1880117;

	wire w740118;
	torch #(1'b1) c740118 (.i_clk(tick), .i_in(), .o_out(w740118));
	wire w780118;
	torch #(1'b1) c780118 (.i_clk(tick), .i_in(), .o_out(w780118));
	wire w820118;
	torch #(1'b1) c820118 (.i_clk(tick), .i_in(), .o_out(w820118));
	wire w860118;
	torch #(1'b1) c860118 (.i_clk(tick), .i_in(), .o_out(w860118));
	wire w900118;
	torch #(1'b1) c900118 (.i_clk(tick), .i_in(), .o_out(w900118));
	wire w940118;
	torch #(1'b1) c940118 (.i_clk(tick), .i_in(), .o_out(w940118));
	wire w980118;
	torch #(1'b1) c980118 (.i_clk(tick), .i_in(), .o_out(w980118));
	wire w1540119;

	wire w1880119;

	wire w1520120;
	repeater #(1, 1'b0, 0, 0) c1520120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520120));
	wire w1640120;
	repeater #(1, 1'b1, 0, 0) c1640120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640120));
	wire w1860120;
	repeater #(1, 1'b1, 0, 0) c1860120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860120));
	wire w1980120;
	repeater #(1, 1'b1, 0, 0) c1980120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980120));
	wire w60121;
	repeater #(2, 1'b0, 0, 0) c60121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60121));
	wire w110121;
	repeater #(2, 1'b0, 0, 0) c110121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110121));
	wire w160121;
	repeater #(2, 1'b0, 0, 0) c160121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160121));
	wire w540121;
	repeater #(2, 1'b0, 0, 0) c540121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540121));
	wire w590121;
	repeater #(2, 1'b1, 0, 0) c590121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590121));
	wire w640121;
	repeater #(2, 1'b1, 0, 0) c640121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640121));
	wire w1430121;
	repeater #(1, 1'b1, 0, 0) c1430121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1430121));
	wire w1590121;
	repeater #(1, 1'b1, 0, 0) c1590121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1590121));
	wire w1770121;
	repeater #(1, 1'b1, 0, 0) c1770121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770121));
	wire w1930121;
	repeater #(1, 1'b1, 0, 0) c1930121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1930121));
	wire w1540122;

	wire w1880122;

	wire w1010123;
	repeater #(1, 1'b0, 0, 0) c1010123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010123));
	wire w1460123;

	wire w1620123;

	wire w1800123;

	wire w1960123;

	wire w1430124;

	wire w1440124;

	wire w1490124;

	wire w1570124;

	wire w1590124;

	wire w1600124;

	wire w1650124;

	wire w1770124;

	wire w1780124;

	wire w1830124;

	wire w1910124;

	wire w1930124;

	wire w1940124;

	wire w1990124;

	wire w710125;
	repeater #(1, 1'b0, 0, 0) c710125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710125));
	wire w1510126;

	wire w1520126;

	wire w1670126;

	wire w1680126;

	wire w1850126;

	wire w1860126;

	wire w2010126;

	wire w2020126;

	wire w260127;
	repeater #(1, 1'b0, 0, 0) c260127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260127));
	wire w440127;
	repeater #(1, 1'b1, 0, 0) c440127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440127));
	wire w800128;
	torch #(1'b1) c800128 (.i_clk(tick), .i_in(), .o_out(w800128));
	wire w840128;
	torch #(1'b1) c840128 (.i_clk(tick), .i_in(), .o_out(w840128));
	wire w880128;
	torch #(1'b1) c880128 (.i_clk(tick), .i_in(), .o_out(w880128));
	wire w920128;
	torch #(1'b1) c920128 (.i_clk(tick), .i_in(), .o_out(w920128));
	wire w1430128;

	wire w1440128;

	wire w1570128;

	wire w1590128;

	wire w1600128;

	wire w1770128;

	wire w1780128;

	wire w1910128;

	wire w1930128;

	wire w1940128;

	wire w330130;
	repeater #(1, 1'b0, 0, 0) c330130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330130));
	wire w1540130;
	torch #(1'b1) c1540130 (.i_clk(tick), .i_in(), .o_out(w1540130));
	wire w1550130;

	wire w1880130;
	torch #(1'b1) c1880130 (.i_clk(tick), .i_in(), .o_out(w1880130));
	wire w1890130;

	wire w80131;
	repeater #(2, 1'b0, 0, 0) c80131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80131));
	wire w620131;
	repeater #(2, 1'b1, 0, 0) c620131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620131));
	wire w1550131;

	wire w1570131;

	wire w1890131;

	wire w1910131;

	wire w50132;
	repeater #(1, 1'b0, 0, 0) c50132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50132));
	wire w130132;
	repeater #(1, 1'b0, 0, 0) c130132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130132));
	wire w140132;
	repeater #(2, 1'b0, 0, 0) c140132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140132));
	wire w370132;

	wire w560132;
	repeater #(2, 1'b0, 0, 0) c560132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560132));
	wire w570132;
	repeater #(1, 1'b0, 0, 0) c570132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570132));
	wire w650132;
	repeater #(1, 1'b1, 0, 0) c650132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650132));
	wire w730132;
	torch #(1'b0) c730132 (.i_clk(tick), .i_in(), .o_out(w730132));
	wire w770132;
	torch #(1'b0) c770132 (.i_clk(tick), .i_in(), .o_out(w770132));
	wire w810132;
	torch #(1'b0) c810132 (.i_clk(tick), .i_in(), .o_out(w810132));
	wire w850132;
	torch #(1'b0) c850132 (.i_clk(tick), .i_in(), .o_out(w850132));
	wire w890132;
	torch #(1'b0) c890132 (.i_clk(tick), .i_in(), .o_out(w890132));
	wire w930132;
	torch #(1'b0) c930132 (.i_clk(tick), .i_in(), .o_out(w930132));
	wire w970132;
	torch #(1'b0) c970132 (.i_clk(tick), .i_in(), .o_out(w970132));
	wire w90133;
	repeater #(1, 1'b0, 0, 0) c90133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90133));
	wire w340133;

	wire w610133;
	repeater #(1, 1'b0, 0, 0) c610133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w610133));
	wire w1570133;

	wire w1580133;

	wire w1590133;

	wire w1910133;

	wire w1920133;

	wire w1930133;

	wire w150134;

	wire w190134;
	repeater #(1, 1'b1, 0, 0) c190134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190134));
	wire w330134;

	wire w350134;
	repeater #(2, 1'b0, 0, 0) c350134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w350134));
	wire w380134;
	repeater #(2, 1'b1, 0, 0) c380134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380134));
	wire w510134;
	repeater #(1, 1'b1, 0, 0) c510134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510134));
	wire w550134;

	wire w740134;
	torch #(1'b1) c740134 (.i_clk(tick), .i_in(), .o_out(w740134));
	wire w780134;
	torch #(1'b1) c780134 (.i_clk(tick), .i_in(), .o_out(w780134));
	wire w820134;
	torch #(1'b1) c820134 (.i_clk(tick), .i_in(), .o_out(w820134));
	wire w860134;
	torch #(1'b1) c860134 (.i_clk(tick), .i_in(), .o_out(w860134));
	wire w900134;
	torch #(1'b1) c900134 (.i_clk(tick), .i_in(), .o_out(w900134));
	wire w940134;
	torch #(1'b1) c940134 (.i_clk(tick), .i_in(), .o_out(w940134));
	wire w980134;
	torch #(1'b1) c980134 (.i_clk(tick), .i_in(), .o_out(w980134));
	wire w1520134;

	wire w1530134;

	wire w1590134;

	wire w1680134;

	wire w1690134;

	wire w1860134;

	wire w1870134;

	wire w1930134;

	wire w2020134;

	wire w2030134;

	wire w160135;

	wire w220135;
	repeater #(2, 1'b0, 0, 0) c220135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220135));
	wire w250135;
	repeater #(2, 1'b0, 0, 0) c250135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250135));
	wire w270135;

	wire w430135;

	wire w450135;
	repeater #(2, 1'b0, 0, 0) c450135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w450135));
	wire w480135;
	repeater #(2, 1'b1, 0, 0) c480135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480135));
	wire w540135;

	wire w150136;
	repeater #(2, 1'b0, 0, 0) c150136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150136));
	wire w260136;

	wire w440136;

	wire w550136;
	repeater #(2, 1'b1, 0, 0) c550136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550136));
	wire w1490136;
	torch #(1'b0) c1490136 (.i_clk(tick), .i_in(), .o_out(w1490136));
	wire w1570136;
	repeater #(1, 1'b1, 0, 0) c1570136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570136));
	wire w1590136;
	torch #(1'b0) c1590136 (.i_clk(tick), .i_in(), .o_out(w1590136));
	wire w1650136;
	torch #(1'b0) c1650136 (.i_clk(tick), .i_in(), .o_out(w1650136));
	wire w1830136;
	torch #(1'b0) c1830136 (.i_clk(tick), .i_in(), .o_out(w1830136));
	wire w1910136;
	repeater #(1, 1'b1, 0, 0) c1910136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910136));
	wire w1930136;
	torch #(1'b0) c1930136 (.i_clk(tick), .i_in(), .o_out(w1930136));
	wire w1990136;
	torch #(1'b0) c1990136 (.i_clk(tick), .i_in(), .o_out(w1990136));
	wire w90137;

	wire w100137;

	wire w230137;

	wire w470137;

	wire w600137;

	wire w610137;

	wire w80138;

	wire w170138;

	wire w530138;

	wire w620138;

	wire w1450138;
	repeater #(1, 1'b1, 0, 0) c1450138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450138));
	wire w1610138;
	repeater #(1, 1'b1, 0, 0) c1610138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610138));
	wire w1790138;
	repeater #(1, 1'b1, 0, 0) c1790138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790138));
	wire w1950138;
	repeater #(1, 1'b1, 0, 0) c1950138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950138));
	wire w410139;
	assign outputs[35] = ();
	wire w1010139;
	repeater #(1, 1'b0, 0, 0) c1010139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010139));
	wire w1580140;
	torch #(1'b1) c1580140 (.i_clk(tick), .i_in(), .o_out(w1580140));
	wire w1920140;
	torch #(1'b1) c1920140 (.i_clk(tick), .i_in(), .o_out(w1920140));
	wire w710141;
	repeater #(1, 1'b0, 0, 0) c710141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710141));
	wire w1500142;
	torch #(1'b1) c1500142 (.i_clk(tick), .i_in(), .o_out(w1500142));
	wire w1660142;
	torch #(1'b1) c1660142 (.i_clk(tick), .i_in(), .o_out(w1660142));
	wire w1840142;
	torch #(1'b1) c1840142 (.i_clk(tick), .i_in(), .o_out(w1840142));
	wire w2000142;
	torch #(1'b1) c2000142 (.i_clk(tick), .i_in(), .o_out(w2000142));
	wire w1570143;
	repeater #(1, 1'b0, 0, 0) c1570143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570143));
	wire w1910143;
	repeater #(1, 1'b0, 0, 0) c1910143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910143));
	wire w800144;
	torch #(1'b1) c800144 (.i_clk(tick), .i_in(), .o_out(w800144));
	wire w840144;
	torch #(1'b1) c840144 (.i_clk(tick), .i_in(), .o_out(w840144));
	wire w880144;
	torch #(1'b1) c880144 (.i_clk(tick), .i_in(), .o_out(w880144));
	wire w920144;
	torch #(1'b1) c920144 (.i_clk(tick), .i_in(), .o_out(w920144));
	wire w1510144;
	repeater #(1, 1'b0, 0, 0) c1510144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510144));
	wire w1670144;
	repeater #(1, 1'b0, 0, 0) c1670144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1670144));
	wire w1850144;
	repeater #(1, 1'b0, 0, 0) c1850144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850144));
	wire w2010144;
	repeater #(1, 1'b0, 0, 0) c2010144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010144));
	wire w1450146;
	repeater #(1, 1'b0, 0, 0) c1450146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450146));
	wire w1790146;
	repeater #(1, 1'b0, 0, 0) c1790146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790146));
	wire w1470147;
	repeater #(1, 1'b0, 0, 0) c1470147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470147));
	wire w1810147;
	repeater #(1, 1'b0, 0, 0) c1810147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810147));
	wire w730148;
	torch #(1'b0) c730148 (.i_clk(tick), .i_in(), .o_out(w730148));
	wire w770148;
	torch #(1'b0) c770148 (.i_clk(tick), .i_in(), .o_out(w770148));
	wire w810148;
	torch #(1'b0) c810148 (.i_clk(tick), .i_in(), .o_out(w810148));
	wire w850148;
	torch #(1'b1) c850148 (.i_clk(tick), .i_in(), .o_out(w850148));
	wire w890148;
	torch #(1'b0) c890148 (.i_clk(tick), .i_in(), .o_out(w890148));
	wire w930148;
	torch #(1'b0) c930148 (.i_clk(tick), .i_in(), .o_out(w930148));
	wire w970148;
	torch #(1'b0) c970148 (.i_clk(tick), .i_in(), .o_out(w970148));
	wire w740150;
	torch #(1'b1) c740150 (.i_clk(tick), .i_in(), .o_out(w740150));
	wire w780150;
	torch #(1'b1) c780150 (.i_clk(tick), .i_in(), .o_out(w780150));
	wire w820150;
	torch #(1'b1) c820150 (.i_clk(tick), .i_in(), .o_out(w820150));
	wire w860150;
	torch #(1'b1) c860150 (.i_clk(tick), .i_in(), .o_out(w860150));
	wire w900150;
	torch #(1'b1) c900150 (.i_clk(tick), .i_in(), .o_out(w900150));
	wire w940150;
	torch #(1'b1) c940150 (.i_clk(tick), .i_in(), .o_out(w940150));
	wire w980150;
	torch #(1'b1) c980150 (.i_clk(tick), .i_in(), .o_out(w980150));
	wire w1010155;
	repeater #(1, 1'b0, 0, 0) c1010155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010155));
	wire w710157;
	repeater #(1, 1'b0, 0, 0) c710157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710157));
	wire w800160;
	torch #(1'b1) c800160 (.i_clk(tick), .i_in(), .o_out(w800160));
	wire w840160;
	torch #(1'b1) c840160 (.i_clk(tick), .i_in(), .o_out(w840160));
	wire w880160;
	torch #(1'b1) c880160 (.i_clk(tick), .i_in(), .o_out(w880160));
	wire w920160;
	torch #(1'b1) c920160 (.i_clk(tick), .i_in(), .o_out(w920160));
	wire w280161;

	wire w460161;

	wire w730164;
	torch #(1'b0) c730164 (.i_clk(tick), .i_in(), .o_out(w730164));
	wire w770164;
	torch #(1'b0) c770164 (.i_clk(tick), .i_in(), .o_out(w770164));
	wire w810164;
	torch #(1'b0) c810164 (.i_clk(tick), .i_in(), .o_out(w810164));
	wire w850164;
	torch #(1'b0) c850164 (.i_clk(tick), .i_in(), .o_out(w850164));
	wire w890164;
	torch #(1'b0) c890164 (.i_clk(tick), .i_in(), .o_out(w890164));
	wire w930164;
	torch #(1'b0) c930164 (.i_clk(tick), .i_in(), .o_out(w930164));
	wire w970164;
	torch #(1'b0) c970164 (.i_clk(tick), .i_in(), .o_out(w970164));
	wire w740166;
	torch #(1'b1) c740166 (.i_clk(tick), .i_in(), .o_out(w740166));
	wire w780166;
	torch #(1'b1) c780166 (.i_clk(tick), .i_in(), .o_out(w780166));
	wire w820166;
	torch #(1'b1) c820166 (.i_clk(tick), .i_in(), .o_out(w820166));
	wire w860166;
	torch #(1'b1) c860166 (.i_clk(tick), .i_in(), .o_out(w860166));
	wire w900166;
	torch #(1'b1) c900166 (.i_clk(tick), .i_in(), .o_out(w900166));
	wire w940166;
	torch #(1'b1) c940166 (.i_clk(tick), .i_in(), .o_out(w940166));
	wire w980166;
	torch #(1'b1) c980166 (.i_clk(tick), .i_in(), .o_out(w980166));
	wire w1010171;
	repeater #(1, 1'b0, 0, 0) c1010171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010171));
	wire w710173;
	repeater #(1, 1'b0, 0, 0) c710173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710173));
	wire w800176;
	torch #(1'b1) c800176 (.i_clk(tick), .i_in(), .o_out(w800176));
	wire w840176;
	torch #(1'b1) c840176 (.i_clk(tick), .i_in(), .o_out(w840176));
	wire w880176;
	torch #(1'b1) c880176 (.i_clk(tick), .i_in(), .o_out(w880176));
	wire w920176;
	torch #(1'b1) c920176 (.i_clk(tick), .i_in(), .o_out(w920176));
	wire w7311;
	torch #(1'b0) c7311 (.i_clk(tick), .i_in(), .o_out(w7311));
	wire w7711;
	torch #(1'b0) c7711 (.i_clk(tick), .i_in(), .o_out(w7711));
	wire w8111;
	torch #(1'b0) c8111 (.i_clk(tick), .i_in(), .o_out(w8111));
	wire w8511;
	torch #(1'b1) c8511 (.i_clk(tick), .i_in(), .o_out(w8511));
	wire w8911;
	torch #(1'b0) c8911 (.i_clk(tick), .i_in(), .o_out(w8911));
	wire w9311;
	torch #(1'b0) c9311 (.i_clk(tick), .i_in(), .o_out(w9311));
	wire w9711;
	torch #(1'b0) c9711 (.i_clk(tick), .i_in(), .o_out(w9711));
	wire w7413;
	torch #(1'b1) c7413 (.i_clk(tick), .i_in(), .o_out(w7413));
	wire w7813;
	torch #(1'b1) c7813 (.i_clk(tick), .i_in(), .o_out(w7813));
	wire w8213;
	torch #(1'b1) c8213 (.i_clk(tick), .i_in(), .o_out(w8213));
	wire w8613;
	torch #(1'b1) c8613 (.i_clk(tick), .i_in(), .o_out(w8613));
	wire w9013;
	torch #(1'b1) c9013 (.i_clk(tick), .i_in(), .o_out(w9013));
	wire w9413;
	torch #(1'b1) c9413 (.i_clk(tick), .i_in(), .o_out(w9413));
	wire w9813;
	torch #(1'b1) c9813 (.i_clk(tick), .i_in(), .o_out(w9813));
	wire w71115;
	repeater #(2, 1'b0, 0, 0) c71115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71115));
	wire w75115;
	repeater #(2, 1'b0, 0, 0) c75115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75115));
	wire w79115;
	repeater #(2, 1'b0, 0, 0) c79115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79115));
	wire w83115;
	repeater #(2, 1'b0, 0, 0) c83115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83115));
	wire w87115;
	repeater #(2, 1'b0, 0, 0) c87115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87115));
	wire w91115;
	repeater #(2, 1'b0, 0, 0) c91115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91115));
	wire w95115;
	repeater #(2, 1'b0, 0, 0) c95115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95115));
	wire w72117;

	wire w76117;

	wire w80117;

	wire w84117;

	wire w88117;

	wire w92117;

	wire w96117;

	wire w72118;

	wire w76118;

	wire w80118;

	wire w84118;

	wire w88118;

	wire w92118;

	wire w96118;

	wire w71121;
	repeater #(1, 1'b1, 0, 0) c71121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71121));
	wire w75121;
	repeater #(1, 1'b1, 0, 0) c75121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75121));
	wire w79121;
	repeater #(1, 1'b1, 0, 0) c79121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79121));
	wire w83121;
	repeater #(1, 1'b1, 0, 0) c83121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83121));
	wire w87121;
	repeater #(1, 1'b1, 0, 0) c87121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87121));
	wire w91121;
	repeater #(1, 1'b1, 0, 0) c91121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91121));
	wire w95121;
	repeater #(1, 1'b1, 0, 0) c95121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95121));
	wire w73122;

	wire w77122;

	wire w81122;

	wire w85122;

	wire w89122;

	wire w93122;

	wire w97122;

	wire w72123;

	wire w76123;

	wire w80123;

	wire w84123;

	wire w88123;

	wire w92123;

	wire w96123;

	wire w74125;
	torch #(1'b1) c74125 (.i_clk(tick), .i_in(), .o_out(w74125));
	wire w78125;
	torch #(1'b0) c78125 (.i_clk(tick), .i_in(), .o_out(w78125));
	wire w82125;
	torch #(1'b0) c82125 (.i_clk(tick), .i_in(), .o_out(w82125));
	wire w86125;
	torch #(1'b1) c86125 (.i_clk(tick), .i_in(), .o_out(w86125));
	wire w90125;
	torch #(1'b0) c90125 (.i_clk(tick), .i_in(), .o_out(w90125));
	wire w94125;
	torch #(1'b0) c94125 (.i_clk(tick), .i_in(), .o_out(w94125));
	wire w98125;
	torch #(1'b0) c98125 (.i_clk(tick), .i_in(), .o_out(w98125));
	wire w99128;
	repeater #(1, 1'b1, 0, 0) c99128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99128));
	wire w100128;
	repeater #(1, 1'b1, 0, 0) c100128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100128));
	wire w84129;
	repeater #(1, 1'b0, 0, 0) c84129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84129));
	wire w99129;
	repeater #(1, 1'b0, 0, 0) c99129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99129));
	wire w74132;

	wire w78132;

	wire w82132;

	wire w86132;

	wire w90132;

	wire w94132;

	wire w98132;

	wire w74134;
	repeater #(1, 1'b0, 0, 0) c74134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74134));
	wire w78134;
	repeater #(1, 1'b0, 0, 0) c78134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78134));
	wire w82134;
	repeater #(1, 1'b0, 0, 0) c82134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82134));
	wire w86134;
	repeater #(1, 1'b0, 0, 0) c86134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86134));
	wire w90134;
	repeater #(1, 1'b0, 0, 0) c90134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90134));
	wire w94134;
	repeater #(1, 1'b0, 0, 0) c94134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94134));
	wire w98134;
	repeater #(1, 1'b0, 0, 0) c98134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98134));
	wire w170163;

	wire w203163;

	wire w204163;

	wire w29164;

	wire w30164;

	wire w63164;

	wire w64164;

	wire w97164;

	wire w171164;
	repeater #(1, 1'b1, 0, 0) c171164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171164));
	wire w205164;
	repeater #(1, 1'b1, 0, 0) c205164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205164));
	wire w31165;
	repeater #(1, 1'b1, 0, 0) c31165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31165));
	wire w65165;
	repeater #(1, 1'b1, 0, 0) c65165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65165));
	wire w168165;

	wire w201165;

	wire w202165;

	wire w27166;

	wire w28166;

	wire w61166;

	wire w62166;

	wire w95166;

	wire w98166;
	repeater #(1, 1'b1, 0, 0) c98166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98166));
	wire w169166;
	repeater #(1, 1'b1, 0, 0) c169166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169166));
	wire w203166;
	repeater #(1, 1'b1, 0, 0) c203166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203166));
	wire w29167;
	repeater #(1, 1'b1, 0, 0) c29167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29167));
	wire w63167;
	repeater #(1, 1'b1, 0, 0) c63167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63167));
	wire w97167;

	wire w166167;

	wire w199167;

	wire w200167;

	wire w25168;

	wire w26168;

	wire w59168;

	wire w60168;

	wire w93168;

	wire w96168;
	repeater #(1, 1'b1, 0, 0) c96168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96168));
	wire w167168;
	repeater #(1, 1'b1, 0, 0) c167168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167168));
	wire w201168;
	repeater #(1, 1'b1, 0, 0) c201168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201168));
	wire w27169;
	repeater #(1, 1'b1, 0, 0) c27169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27169));
	wire w61169;
	repeater #(1, 1'b1, 0, 0) c61169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61169));
	wire w95169;

	wire w164169;

	wire w197169;

	wire w198169;

	wire w23170;

	wire w24170;

	wire w57170;

	wire w58170;

	wire w91170;

	wire w94170;
	repeater #(1, 1'b1, 0, 0) c94170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94170));
	wire w165170;
	repeater #(1, 1'b1, 0, 0) c165170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165170));
	wire w199170;
	repeater #(1, 1'b1, 0, 0) c199170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199170));
	wire w25171;
	repeater #(1, 1'b1, 0, 0) c25171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25171));
	wire w59171;
	repeater #(1, 1'b1, 0, 0) c59171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59171));
	wire w93171;

	wire w162171;

	wire w195171;

	wire w196171;

	wire w21172;

	wire w22172;

	wire w55172;

	wire w56172;

	wire w89172;

	wire w92172;
	repeater #(1, 1'b1, 0, 0) c92172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92172));
	wire w163172;
	repeater #(1, 1'b1, 0, 0) c163172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163172));
	wire w197172;
	repeater #(1, 1'b1, 0, 0) c197172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197172));
	wire w23173;
	repeater #(1, 1'b1, 0, 0) c23173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23173));
	wire w57173;
	repeater #(1, 1'b1, 0, 0) c57173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57173));
	wire w91173;

	wire w160173;

	wire w193173;

	wire w194173;

	wire w19174;

	wire w20174;

	wire w53174;

	wire w54174;

	wire w87174;

	wire w90174;
	repeater #(1, 1'b1, 0, 0) c90174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90174));
	wire w161174;
	repeater #(1, 1'b1, 0, 0) c161174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161174));
	wire w195174;
	repeater #(1, 1'b1, 0, 0) c195174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195174));
	wire w21175;
	repeater #(1, 1'b1, 0, 0) c21175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21175));
	wire w55175;
	repeater #(1, 1'b1, 0, 0) c55175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55175));
	wire w89175;

	wire w158175;

	wire w191175;

	wire w192175;

	wire w17176;

	wire w18176;

	wire w51176;

	wire w52176;

	wire w85176;

	wire w88176;
	repeater #(1, 1'b1, 0, 0) c88176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88176));
	wire w159176;
	repeater #(1, 1'b1, 0, 0) c159176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159176));
	wire w193176;
	repeater #(1, 1'b1, 0, 0) c193176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193176));
	wire w19177;
	repeater #(1, 1'b1, 0, 0) c19177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19177));
	wire w53177;
	repeater #(1, 1'b1, 0, 0) c53177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53177));
	wire w87177;

	wire w156177;

	wire w189177;

	wire w190177;

	wire w15178;

	wire w16178;

	wire w49178;

	wire w50178;

	wire w83178;

	wire w86178;
	repeater #(1, 1'b1, 0, 0) c86178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86178));
	wire w157178;
	repeater #(1, 1'b0, 0, 0) c157178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157178));
	wire w191178;
	repeater #(1, 1'b0, 0, 0) c191178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191178));
	wire w17179;
	repeater #(1, 1'b0, 0, 0) c17179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17179));
	wire w51179;
	repeater #(1, 1'b0, 0, 0) c51179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51179));
	wire w85179;

	wire w154179;

	wire w187179;

	wire w188179;

	wire w13180;

	wire w14180;

	wire w47180;

	wire w48180;

	wire w81180;

	wire w84180;
	repeater #(1, 1'b0, 0, 0) c84180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84180));
	wire w155180;
	repeater #(1, 1'b1, 0, 0) c155180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155180));
	wire w189180;
	repeater #(1, 1'b1, 0, 0) c189180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189180));
	wire w15181;
	repeater #(1, 1'b1, 0, 0) c15181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15181));
	wire w49181;
	repeater #(1, 1'b1, 0, 0) c49181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49181));
	wire w83181;

	wire w152181;

	wire w185181;

	wire w186181;

	wire w11182;

	wire w12182;

	wire w45182;

	wire w46182;

	wire w79182;

	wire w82182;
	repeater #(1, 1'b1, 0, 0) c82182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82182));
	wire w153182;
	repeater #(1, 1'b1, 0, 0) c153182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153182));
	wire w187182;
	repeater #(1, 1'b1, 0, 0) c187182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187182));
	wire w13183;
	repeater #(1, 1'b1, 0, 0) c13183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13183));
	wire w47183;
	repeater #(1, 1'b1, 0, 0) c47183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47183));
	wire w81183;

	wire w150183;

	wire w183183;

	wire w184183;

	wire w9184;

	wire w10184;

	wire w43184;

	wire w44184;

	wire w77184;

	wire w80184;
	repeater #(1, 1'b1, 0, 0) c80184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80184));
	wire w151184;
	repeater #(1, 1'b1, 0, 0) c151184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151184));
	wire w185184;
	repeater #(1, 1'b1, 0, 0) c185184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185184));
	wire w11185;
	repeater #(1, 1'b1, 0, 0) c11185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11185));
	wire w45185;
	repeater #(1, 1'b1, 0, 0) c45185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45185));
	wire w79185;

	wire w148185;

	wire w181185;

	wire w182185;

	wire w7186;

	wire w8186;

	wire w41186;

	wire w42186;

	wire w75186;

	wire w78186;
	repeater #(1, 1'b1, 0, 0) c78186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78186));
	wire w149186;
	repeater #(1, 1'b1, 0, 0) c149186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149186));
	wire w183186;
	repeater #(1, 1'b1, 0, 0) c183186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183186));
	wire w9187;
	repeater #(1, 1'b1, 0, 0) c9187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9187));
	wire w43187;
	repeater #(1, 1'b1, 0, 0) c43187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43187));
	wire w77187;

	wire w146187;

	wire w179187;

	wire w180187;

	wire w5188;

	wire w6188;

	wire w39188;

	wire w40188;

	wire w73188;

	wire w76188;
	repeater #(1, 1'b1, 0, 0) c76188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76188));
	wire w147188;
	repeater #(1, 1'b1, 0, 0) c147188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147188));
	wire w181188;
	repeater #(1, 1'b1, 0, 0) c181188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181188));
	wire w7189;
	repeater #(1, 1'b1, 0, 0) c7189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7189));
	wire w41189;
	repeater #(1, 1'b1, 0, 0) c41189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41189));
	wire w75189;

	wire w177189;

	wire w3190;

	wire w37190;

	wire w71190;

	wire w74190;
	repeater #(1, 1'b1, 0, 0) c74190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74190));
	wire w145190;
	repeater #(1, 1'b1, 0, 0) c145190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145190));
	wire w179190;
	repeater #(1, 1'b1, 0, 0) c179190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179190));
	wire w5191;
	repeater #(1, 1'b1, 0, 0) c5191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5191));
	wire w39191;
	repeater #(1, 1'b1, 0, 0) c39191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39191));
	wire w73191;

	wire w72192;
	repeater #(2, 1'b1, 0, 0) c72192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72192));
	wire w74193;
	repeater #(1, 1'b1, 0, 0) c74193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74193));
	wire w164195;
	repeater #(2, 1'b1, 0, 0) c164195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164195));
	wire w198195;
	repeater #(2, 1'b1, 0, 0) c198195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198195));
	wire w73196;
	torch #(1'b1) c73196 (.i_clk(tick), .i_in(), .o_out(w73196));
	wire w77196;
	torch #(1'b1) c77196 (.i_clk(tick), .i_in(), .o_out(w77196));
	wire w81196;
	torch #(1'b1) c81196 (.i_clk(tick), .i_in(), .o_out(w81196));
	wire w85196;
	torch #(1'b0) c85196 (.i_clk(tick), .i_in(), .o_out(w85196));
	wire w89196;
	torch #(1'b1) c89196 (.i_clk(tick), .i_in(), .o_out(w89196));
	wire w93196;
	torch #(1'b1) c93196 (.i_clk(tick), .i_in(), .o_out(w93196));
	wire w97196;
	torch #(1'b1) c97196 (.i_clk(tick), .i_in(), .o_out(w97196));
	wire w150197;
	repeater #(1, 1'b1, 0, 0) c150197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150197));
	wire w156197;
	torch #(1'b0) c156197 (.i_clk(tick), .i_in(), .o_out(w156197));
	wire w166197;
	repeater #(1, 1'b1, 0, 0) c166197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166197));
	wire w184197;
	repeater #(1, 1'b1, 0, 0) c184197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184197));
	wire w190197;
	torch #(1'b0) c190197 (.i_clk(tick), .i_in(), .o_out(w190197));
	wire w200197;
	repeater #(1, 1'b1, 0, 0) c200197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200197));
	wire w74199;
	repeater #(1, 1'b1, 0, 0) c74199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74199));
	wire w78199;
	repeater #(1, 1'b1, 0, 0) c78199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78199));
	wire w82199;
	repeater #(1, 1'b1, 0, 0) c82199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82199));
	wire w86199;
	repeater #(1, 1'b0, 0, 0) c86199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86199));
	wire w90199;
	repeater #(1, 1'b1, 0, 0) c90199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90199));
	wire w94199;
	repeater #(1, 1'b1, 0, 0) c94199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94199));
	wire w98199;
	repeater #(1, 1'b1, 0, 0) c98199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98199));
	wire w731100;
	torch #(1'b1) c731100 (.i_clk(tick), .i_in(), .o_out(w731100));
	wire w771100;
	torch #(1'b1) c771100 (.i_clk(tick), .i_in(), .o_out(w771100));
	wire w811100;
	torch #(1'b1) c811100 (.i_clk(tick), .i_in(), .o_out(w811100));
	wire w851100;
	torch #(1'b0) c851100 (.i_clk(tick), .i_in(), .o_out(w851100));
	wire w891100;
	torch #(1'b1) c891100 (.i_clk(tick), .i_in(), .o_out(w891100));
	wire w931100;
	torch #(1'b1) c931100 (.i_clk(tick), .i_in(), .o_out(w931100));
	wire w971100;
	torch #(1'b1) c971100 (.i_clk(tick), .i_in(), .o_out(w971100));
	wire w1451100;
	repeater #(1, 1'b1, 0, 0) c1451100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1451100));
	wire w1571100;
	repeater #(1, 1'b0, 0, 0) c1571100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1571100));
	wire w1791100;
	repeater #(1, 1'b1, 0, 0) c1791100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1791100));
	wire w1911100;
	repeater #(1, 1'b1, 0, 0) c1911100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911100));
	wire w1501101;
	repeater #(1, 1'b1, 0, 0) c1501101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1501101));
	wire w1661101;
	repeater #(1, 1'b1, 0, 0) c1661101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661101));
	wire w1841101;
	repeater #(1, 1'b1, 0, 0) c1841101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1841101));
	wire w2001101;
	repeater #(1, 1'b1, 0, 0) c2001101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2001101));
	wire w111102;
	torch #(1'b0) c111102 (.i_clk(tick), .i_in(), .o_out(w111102));
	wire w151102;
	torch #(1'b1) c151102 (.i_clk(tick), .i_in(), .o_out(w151102));
	wire w191102;
	torch #(1'b1) c191102 (.i_clk(tick), .i_in(), .o_out(w191102));
	wire w231102;
	torch #(1'b0) c231102 (.i_clk(tick), .i_in(), .o_out(w231102));
	wire w471102;
	torch #(1'b0) c471102 (.i_clk(tick), .i_in(), .o_out(w471102));
	wire w511102;
	torch #(1'b0) c511102 (.i_clk(tick), .i_in(), .o_out(w511102));
	wire w551102;
	torch #(1'b0) c551102 (.i_clk(tick), .i_in(), .o_out(w551102));
	wire w591102;
	torch #(1'b1) c591102 (.i_clk(tick), .i_in(), .o_out(w591102));
	wire w1551102;

	wire w1891102;

	wire w721103;
	torch #(1'b0) c721103 (.i_clk(tick), .i_in(), .o_out(w721103));
	wire w761103;
	torch #(1'b0) c761103 (.i_clk(tick), .i_in(), .o_out(w761103));
	wire w801103;
	torch #(1'b0) c801103 (.i_clk(tick), .i_in(), .o_out(w801103));
	wire w841103;
	torch #(1'b1) c841103 (.i_clk(tick), .i_in(), .o_out(w841103));
	wire w881103;
	torch #(1'b0) c881103 (.i_clk(tick), .i_in(), .o_out(w881103));
	wire w921103;
	torch #(1'b0) c921103 (.i_clk(tick), .i_in(), .o_out(w921103));
	wire w961103;
	torch #(1'b0) c961103 (.i_clk(tick), .i_in(), .o_out(w961103));
	wire w1471103;

	wire w1631103;

	wire w1811103;

	wire w1971103;

	wire w1441104;

	wire w1491104;

	wire w1501104;

	wire w1601104;

	wire w1651104;

	wire w1661104;

	wire w1781104;

	wire w1831104;

	wire w1841104;

	wire w1941104;

	wire w1991104;

	wire w2001104;

	wire w1421106;

	wire w1581106;

	wire w1761106;

	wire w1921106;

	wire w1481107;

	wire w1491107;

	wire w1641107;

	wire w1651107;

	wire w1821107;

	wire w1831107;

	wire w1981107;

	wire w1991107;

	wire w1581108;

	wire w1921108;

	wire w111109;
	repeater #(2, 1'b1, 0, 0) c111109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111109));
	wire w131109;
	repeater #(1, 1'b0, 0, 0) c131109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131109));
	wire w151109;
	repeater #(2, 1'b0, 0, 0) c151109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151109));
	wire w171109;
	repeater #(1, 1'b0, 0, 0) c171109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171109));
	wire w191109;
	repeater #(2, 1'b0, 0, 0) c191109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191109));
	wire w211109;
	repeater #(1, 1'b0, 0, 0) c211109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w211109));
	wire w231109;
	repeater #(2, 1'b1, 0, 0) c231109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w231109));
	wire w251109;
	repeater #(1, 1'b0, 0, 0) c251109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w251109));
	wire w451109;
	repeater #(1, 1'b1, 0, 0) c451109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w451109));
	wire w471109;
	repeater #(2, 1'b1, 0, 0) c471109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w471109));
	wire w491109;
	repeater #(1, 1'b1, 0, 0) c491109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w491109));
	wire w511109;
	repeater #(2, 1'b1, 0, 0) c511109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w511109));
	wire w531109;
	repeater #(1, 1'b1, 0, 0) c531109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w531109));
	wire w551109;
	repeater #(2, 1'b1, 0, 0) c551109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w551109));
	wire w571109;
	repeater #(1, 1'b1, 0, 0) c571109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w571109));
	wire w591109;
	repeater #(2, 1'b0, 0, 0) c591109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w591109));
	wire w801109;
	torch #(1'b1) c801109 (.i_clk(tick), .i_in(), .o_out(w801109));
	wire w841109;
	torch #(1'b1) c841109 (.i_clk(tick), .i_in(), .o_out(w841109));
	wire w881109;
	torch #(1'b1) c881109 (.i_clk(tick), .i_in(), .o_out(w881109));
	wire w921109;
	torch #(1'b1) c921109 (.i_clk(tick), .i_in(), .o_out(w921109));
	wire w1421110;

	wire w1461110;

	wire w1501110;

	wire w1541110;

	wire w1581110;

	wire w1621110;

	wire w1661110;

	wire w1761110;

	wire w1801110;

	wire w1841110;

	wire w1881110;

	wire w1921110;

	wire w1961110;

	wire w2001110;

	wire w201111;

	wire w501111;

	wire w121112;

	wire w161112;

	wire w191112;

	wire w211112;

	wire w241112;

	wire w461112;

	wire w491112;

	wire w511112;

	wire w541112;

	wire w581112;

	wire w111113;

	wire w131113;

	wire w151113;

	wire w171113;

	wire w201113;

	wire w231113;

	wire w251113;

	wire w451113;

	wire w471113;

	wire w501113;

	wire w531113;

	wire w551113;

	wire w571113;

	wire w591113;

	wire w161114;

	wire w541114;

	wire w1421114;

	wire w1461114;

	wire w1501114;

	wire w1541114;

	wire w1581114;

	wire w1621114;

	wire w1661114;

	wire w1761114;

	wire w1801114;

	wire w1841114;

	wire w1881114;

	wire w1921114;

	wire w1961114;

	wire w2001114;

	wire w121115;

	wire w161115;

	wire w171115;

	wire w211115;

	wire w231115;

	wire w251115;

	wire w451115;

	wire w471115;

	wire w491115;

	wire w531115;

	wire w541115;

	wire w581115;

	wire w161116;

	wire w541116;

	wire w1401116;
	repeater #(1, 1'b1, 0, 0) c1401116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401116));
	wire w1441116;
	repeater #(1, 1'b1, 0, 0) c1441116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441116));
	wire w1481116;
	repeater #(1, 1'b1, 0, 0) c1481116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1481116));
	wire w1521116;
	repeater #(1, 1'b0, 0, 0) c1521116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1521116));
	wire w1741116;
	repeater #(1, 1'b1, 0, 0) c1741116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741116));
	wire w1781116;
	repeater #(1, 1'b1, 0, 0) c1781116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781116));
	wire w1821116;
	repeater #(1, 1'b1, 0, 0) c1821116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821116));
	wire w1861116;
	repeater #(1, 1'b1, 0, 0) c1861116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861116));
	wire w131117;

	wire w151117;

	wire w551117;

	wire w571117;

	wire w1581117;

	wire w1621117;

	wire w1661117;

	wire w1921117;

	wire w1961117;

	wire w2001117;

	wire w731118;
	torch #(1'b1) c731118 (.i_clk(tick), .i_in(), .o_out(w731118));
	wire w771118;
	torch #(1'b1) c771118 (.i_clk(tick), .i_in(), .o_out(w771118));
	wire w811118;
	torch #(1'b1) c811118 (.i_clk(tick), .i_in(), .o_out(w811118));
	wire w851118;
	torch #(1'b0) c851118 (.i_clk(tick), .i_in(), .o_out(w851118));
	wire w891118;
	torch #(1'b1) c891118 (.i_clk(tick), .i_in(), .o_out(w891118));
	wire w931118;
	torch #(1'b1) c931118 (.i_clk(tick), .i_in(), .o_out(w931118));
	wire w971118;
	torch #(1'b1) c971118 (.i_clk(tick), .i_in(), .o_out(w971118));
	wire w741119;
	repeater #(1, 1'b0, 0, 0) c741119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741119));
	wire w781119;
	repeater #(1, 1'b0, 0, 0) c781119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w781119));
	wire w821119;
	repeater #(1, 1'b0, 0, 0) c821119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821119));
	wire w861119;
	repeater #(1, 1'b1, 0, 0) c861119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861119));
	wire w901119;
	repeater #(1, 1'b0, 0, 0) c901119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901119));
	wire w941119;
	repeater #(1, 1'b0, 0, 0) c941119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941119));
	wire w981119;
	repeater #(1, 1'b0, 0, 0) c981119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981119));
	wire w1581119;

	wire w1921119;

	wire w1401120;
	repeater #(1, 1'b1, 0, 0) c1401120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401120));
	wire w1561120;
	repeater #(1, 1'b1, 0, 0) c1561120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1561120));
	wire w1741120;
	repeater #(1, 1'b1, 0, 0) c1741120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741120));
	wire w1901120;
	repeater #(1, 1'b1, 0, 0) c1901120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901120));
	wire w721121;

	wire w741121;
	repeater #(1, 1'b0, 0, 0) c741121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741121));
	wire w761121;

	wire w781121;
	repeater #(1, 1'b0, 0, 0) c781121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w781121));
	wire w801121;

	wire w821121;
	repeater #(1, 1'b0, 0, 0) c821121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821121));
	wire w841121;

	wire w861121;
	repeater #(1, 1'b1, 0, 0) c861121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861121));
	wire w881121;

	wire w901121;
	repeater #(1, 1'b0, 0, 0) c901121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901121));
	wire w921121;

	wire w941121;
	repeater #(1, 1'b0, 0, 0) c941121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941121));
	wire w961121;

	wire w981121;
	repeater #(1, 1'b0, 0, 0) c981121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981121));
	wire w1471121;
	repeater #(1, 1'b1, 0, 0) c1471121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1471121));
	wire w1631121;
	repeater #(1, 1'b1, 0, 0) c1631121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1631121));
	wire w1811121;
	repeater #(1, 1'b1, 0, 0) c1811121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1811121));
	wire w1971121;
	repeater #(1, 1'b1, 0, 0) c1971121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1971121));
	wire w1421122;

	wire w1581122;

	wire w1761122;

	wire w1921122;

	wire w1501123;

	wire w1841123;

	wire w1451124;

	wire w1471124;

	wire w1481124;

	wire w1531124;

	wire w1611124;

	wire w1631124;

	wire w1641124;

	wire w1791124;

	wire w1811124;

	wire w1821124;

	wire w1871124;

	wire w1951124;

	wire w1971124;

	wire w1981124;

	wire w801125;
	torch #(1'b1) c801125 (.i_clk(tick), .i_in(), .o_out(w801125));
	wire w841125;
	torch #(1'b1) c841125 (.i_clk(tick), .i_in(), .o_out(w841125));
	wire w881125;
	torch #(1'b1) c881125 (.i_clk(tick), .i_in(), .o_out(w881125));
	wire w921125;
	torch #(1'b1) c921125 (.i_clk(tick), .i_in(), .o_out(w921125));
	wire w1551126;

	wire w1561126;

	wire w1891126;

	wire w1901126;

	wire w1451128;

	wire w1471128;

	wire w1481128;

	wire w1611128;

	wire w1631128;

	wire w1641128;

	wire w1791128;

	wire w1811128;

	wire w1821128;

	wire w1951128;

	wire w1971128;

	wire w1981128;

	wire w241130;
	repeater #(1, 1'b0, 0, 0) c241130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w241130));
	wire w461130;
	repeater #(1, 1'b1, 0, 0) c461130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w461130));
	wire w1421130;
	torch #(1'b1) c1421130 (.i_clk(tick), .i_in(), .o_out(w1421130));
	wire w1431130;

	wire w1581130;
	torch #(1'b1) c1581130 (.i_clk(tick), .i_in(), .o_out(w1581130));
	wire w1591130;

	wire w1761130;
	torch #(1'b1) c1761130 (.i_clk(tick), .i_in(), .o_out(w1761130));
	wire w1771130;

	wire w1921130;
	torch #(1'b1) c1921130 (.i_clk(tick), .i_in(), .o_out(w1921130));
	wire w1931130;

	wire w351131;

	wire w1431131;

	wire w1451131;

	wire w1591131;

	wire w1611131;

	wire w1771131;

	wire w1791131;

	wire w1931131;

	wire w1951131;

	wire w361132;

	wire w131133;

	wire w271133;
	repeater #(1, 1'b0, 0, 0) c271133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w271133));
	wire w281133;

	wire w361133;
	repeater #(1, 1'b0, 0, 0) c361133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w361133));
	wire w421133;

	wire w431133;
	repeater #(1, 1'b0, 0, 0) c431133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w431133));
	wire w571133;

	wire w1451133;

	wire w1461133;

	wire w1471133;

	wire w1611133;

	wire w1621133;

	wire w1631133;

	wire w1791133;

	wire w1801133;

	wire w1811133;

	wire w1951133;

	wire w1961133;

	wire w1971133;

	wire w131134;
	repeater #(1, 1'b0, 0, 0) c131134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131134));
	wire w241134;

	wire w251134;

	wire w451134;

	wire w461134;

	wire w571134;
	repeater #(1, 1'b1, 0, 0) c571134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w571134));
	wire w731134;
	torch #(1'b1) c731134 (.i_clk(tick), .i_in(), .o_out(w731134));
	wire w771134;
	torch #(1'b1) c771134 (.i_clk(tick), .i_in(), .o_out(w771134));
	wire w811134;
	torch #(1'b1) c811134 (.i_clk(tick), .i_in(), .o_out(w811134));
	wire w851134;
	torch #(1'b1) c851134 (.i_clk(tick), .i_in(), .o_out(w851134));
	wire w891134;
	torch #(1'b1) c891134 (.i_clk(tick), .i_in(), .o_out(w891134));
	wire w931134;
	torch #(1'b1) c931134 (.i_clk(tick), .i_in(), .o_out(w931134));
	wire w971134;
	torch #(1'b1) c971134 (.i_clk(tick), .i_in(), .o_out(w971134));
	wire w1471134;

	wire w1561134;

	wire w1571134;

	wire w1631134;

	wire w1811134;

	wire w1901134;

	wire w1911134;

	wire w1971134;

	wire w351135;

	wire w361135;

	wire w741135;
	repeater #(1, 1'b0, 0, 0) c741135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741135));
	wire w781135;
	repeater #(1, 1'b0, 0, 0) c781135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w781135));
	wire w821135;
	repeater #(1, 1'b0, 0, 0) c821135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821135));
	wire w861135;
	repeater #(1, 1'b1, 0, 0) c861135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861135));
	wire w901135;
	repeater #(1, 1'b0, 0, 0) c901135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901135));
	wire w941135;
	repeater #(1, 1'b0, 0, 0) c941135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941135));
	wire w981135;
	repeater #(1, 1'b0, 0, 0) c981135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981135));
	wire w141136;

	wire w200;

	wire w800;
	repeater #(1, 1'b0, 0, 0) c800 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800));
	wire w1600;

	wire w1700;
	repeater #(1, 1'b0, 0, 0) c1700 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1700));
	wire w3000;
	repeater #(1, 1'b0, 0, 0) c3000 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3000));
	wire w3600;

	wire w4000;

	wire w12900;
	repeater #(1, 1'b0, 0, 0) c12900 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12900));
	wire w13100;
	torch #(1'b0) c13100 (.i_clk(tick), .i_in(), .o_out(w13100));
	wire w13700;
	torch #(1'b0) c13700 (.i_clk(tick), .i_in(), .o_out(w13700));
	wire w14500;
	repeater #(1, 1'b0, 0, 0) c14500 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14500));
	wire w14700;
	torch #(1'b0) c14700 (.i_clk(tick), .i_in(), .o_out(w14700));
	wire w15300;
	torch #(1'b0) c15300 (.i_clk(tick), .i_in(), .o_out(w15300));
	wire w16300;
	repeater #(1, 1'b0, 0, 0) c16300 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16300));
	wire w16500;
	torch #(1'b0) c16500 (.i_clk(tick), .i_in(), .o_out(w16500));
	wire w17100;
	torch #(1'b0) c17100 (.i_clk(tick), .i_in(), .o_out(w17100));
	wire w17900;
	repeater #(1, 1'b0, 0, 0) c17900 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17900));
	wire w18100;
	torch #(1'b0) c18100 (.i_clk(tick), .i_in(), .o_out(w18100));
	wire w18700;
	torch #(1'b0) c18700 (.i_clk(tick), .i_in(), .o_out(w18700));
	wire w20600;

	wire w001;
	repeater #(1, 1'b0, 0, 0) c001 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w001));
	wire w101;

	wire w801;

	wire w2501;

	wire w3001;

	wire w3701;

	wire w3801;
	repeater #(1, 1'b1, 0, 0) c3801 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3801));
	wire w4001;

	wire w5601;

	wire w5801;
	repeater #(1, 1'b0, 0, 0) c5801 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5801));
	wire w6001;

	wire w6201;
	repeater #(1, 1'b0, 0, 0) c6201 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6201));
	wire w6401;

	wire w6601;
	repeater #(1, 1'b0, 0, 0) c6601 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6601));
	wire w6801;

	wire w7001;
	repeater #(1, 1'b1, 0, 0) c7001 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7001));
	wire w7201;

	wire w7401;
	repeater #(1, 1'b0, 0, 0) c7401 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7401));
	wire w7601;

	wire w7801;
	repeater #(1, 1'b0, 0, 0) c7801 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7801));
	wire w8001;

	wire w8201;
	repeater #(1, 1'b0, 0, 0) c8201 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8201));
	wire w902;

	wire w1302;
	repeater #(1, 1'b0, 0, 0) c1302 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1302));
	wire w2602;
	repeater #(2, 1'b1, 0, 0) c2602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2602));
	wire w2902;

	wire w13302;
	repeater #(1, 1'b1, 0, 0) c13302 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13302));
	wire w14902;
	repeater #(1, 1'b1, 0, 0) c14902 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14902));
	wire w16702;
	repeater #(1, 1'b1, 0, 0) c16702 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16702));
	wire w18302;
	repeater #(1, 1'b1, 0, 0) c18302 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18302));
	wire w1203;
	assign outputs[36] = ();
	wire w13004;
	torch #(1'b1) c13004 (.i_clk(tick), .i_in(), .o_out(w13004));
	wire w14604;
	torch #(1'b1) c14604 (.i_clk(tick), .i_in(), .o_out(w14604));
	wire w16404;
	torch #(1'b1) c16404 (.i_clk(tick), .i_in(), .o_out(w16404));
	wire w18004;
	torch #(1'b1) c18004 (.i_clk(tick), .i_in(), .o_out(w18004));
	wire w6405;
	torch #(1'b1) c6405 (.i_clk(tick), .i_in(), .o_out(w6405));
	wire w6805;
	torch #(1'b1) c6805 (.i_clk(tick), .i_in(), .o_out(w6805));
	wire w7205;
	torch #(1'b1) c7205 (.i_clk(tick), .i_in(), .o_out(w7205));
	wire w7605;
	torch #(1'b1) c7605 (.i_clk(tick), .i_in(), .o_out(w7605));
	wire w13806;
	torch #(1'b1) c13806 (.i_clk(tick), .i_in(), .o_out(w13806));
	wire w15406;
	torch #(1'b1) c15406 (.i_clk(tick), .i_in(), .o_out(w15406));
	wire w17206;
	torch #(1'b1) c17206 (.i_clk(tick), .i_in(), .o_out(w17206));
	wire w18806;
	torch #(1'b1) c18806 (.i_clk(tick), .i_in(), .o_out(w18806));
	wire w12907;
	repeater #(2, 1'b0, 0, 0) c12907 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12907));
	wire w14507;
	repeater #(1, 1'b0, 0, 0) c14507 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14507));
	wire w16307;
	repeater #(2, 1'b0, 0, 0) c16307 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16307));
	wire w17907;
	repeater #(1, 1'b0, 0, 0) c17907 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17907));
	wire w13908;
	repeater #(1, 1'b0, 0, 0) c13908 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13908));
	wire w15508;
	repeater #(1, 1'b0, 0, 0) c15508 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15508));
	wire w17308;
	repeater #(1, 1'b0, 0, 0) c17308 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17308));
	wire w18908;
	repeater #(1, 1'b0, 0, 0) c18908 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18908));
	wire w133010;
	repeater #(1, 1'b0, 0, 0) c133010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133010));
	wire w167010;
	repeater #(1, 1'b0, 0, 0) c167010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167010));
	wire w135011;
	repeater #(1, 1'b0, 0, 0) c135011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135011));
	wire w169011;
	repeater #(1, 1'b0, 0, 0) c169011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169011));
	wire w57014;
	torch #(1'b1) c57014 (.i_clk(tick), .i_in(), .o_out(w57014));
	wire w61014;
	torch #(1'b1) c61014 (.i_clk(tick), .i_in(), .o_out(w61014));
	wire w65014;
	torch #(1'b1) c65014 (.i_clk(tick), .i_in(), .o_out(w65014));
	wire w69014;
	torch #(1'b0) c69014 (.i_clk(tick), .i_in(), .o_out(w69014));
	wire w73014;
	torch #(1'b1) c73014 (.i_clk(tick), .i_in(), .o_out(w73014));
	wire w77014;
	torch #(1'b1) c77014 (.i_clk(tick), .i_in(), .o_out(w77014));
	wire w81014;
	torch #(1'b1) c81014 (.i_clk(tick), .i_in(), .o_out(w81014));
	wire w58015;
	repeater #(1, 1'b0, 0, 0) c58015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58015));
	wire w62015;
	repeater #(1, 1'b0, 0, 0) c62015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62015));
	wire w66015;
	repeater #(1, 1'b0, 0, 0) c66015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66015));
	wire w70015;
	repeater #(1, 1'b1, 0, 0) c70015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70015));
	wire w74015;
	repeater #(1, 1'b0, 0, 0) c74015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74015));
	wire w78015;
	repeater #(1, 1'b0, 0, 0) c78015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78015));
	wire w82015;
	repeater #(1, 1'b0, 0, 0) c82015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82015));
	wire w56017;

	wire w58017;
	repeater #(1, 1'b0, 0, 0) c58017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58017));
	wire w60017;

	wire w62017;
	repeater #(1, 1'b0, 0, 0) c62017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62017));
	wire w64017;

	wire w66017;
	repeater #(1, 1'b0, 0, 0) c66017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66017));
	wire w68017;

	wire w70017;
	repeater #(1, 1'b1, 0, 0) c70017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70017));
	wire w72017;

	wire w74017;
	repeater #(1, 1'b0, 0, 0) c74017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74017));
	wire w76017;

	wire w78017;
	repeater #(1, 1'b0, 0, 0) c78017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78017));
	wire w80017;

	wire w82017;
	repeater #(1, 1'b0, 0, 0) c82017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82017));
	wire w64021;
	torch #(1'b1) c64021 (.i_clk(tick), .i_in(), .o_out(w64021));
	wire w68021;
	torch #(1'b1) c68021 (.i_clk(tick), .i_in(), .o_out(w68021));
	wire w72021;
	torch #(1'b1) c72021 (.i_clk(tick), .i_in(), .o_out(w72021));
	wire w76021;
	torch #(1'b1) c76021 (.i_clk(tick), .i_in(), .o_out(w76021));
	wire w18025;

	wire w19025;
	repeater #(1, 1'b0, 0, 0) c19025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19025));
	wire w20026;
	repeater #(1, 1'b0, 0, 0) c20026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20026));
	wire w23026;
	repeater #(2, 1'b0, 0, 0) c23026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23026));
	wire w15027;
	repeater #(1, 1'b0, 0, 0) c15027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15027));
	wire w28027;
	repeater #(2, 1'b0, 0, 0) c28027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28027));
	wire w14028;
	assign outputs[37] = ();
	wire w17028;

	wire w26028;

	wire w17029;

	wire w26029;

	wire w15030;
	repeater #(1, 1'b0, 0, 0) c15030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15030));
	wire w28030;
	repeater #(1, 1'b0, 0, 0) c28030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28030));
	wire w57030;
	torch #(1'b1) c57030 (.i_clk(tick), .i_in(), .o_out(w57030));
	wire w61030;
	torch #(1'b1) c61030 (.i_clk(tick), .i_in(), .o_out(w61030));
	wire w65030;
	torch #(1'b1) c65030 (.i_clk(tick), .i_in(), .o_out(w65030));
	wire w69030;
	torch #(1'b1) c69030 (.i_clk(tick), .i_in(), .o_out(w69030));
	wire w73030;
	torch #(1'b1) c73030 (.i_clk(tick), .i_in(), .o_out(w73030));
	wire w77030;
	torch #(1'b1) c77030 (.i_clk(tick), .i_in(), .o_out(w77030));
	wire w81030;
	torch #(1'b1) c81030 (.i_clk(tick), .i_in(), .o_out(w81030));
	wire w58031;
	repeater #(1, 1'b0, 0, 0) c58031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58031));
	wire w62031;
	repeater #(1, 1'b0, 0, 0) c62031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62031));
	wire w66031;
	repeater #(1, 1'b0, 0, 0) c66031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66031));
	wire w70031;
	repeater #(1, 1'b1, 0, 0) c70031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70031));
	wire w74031;
	repeater #(1, 1'b0, 0, 0) c74031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74031));
	wire w78031;
	repeater #(1, 1'b0, 0, 0) c78031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78031));
	wire w82031;
	repeater #(1, 1'b0, 0, 0) c82031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82031));
	wire w56033;

	wire w58033;
	repeater #(1, 1'b0, 0, 0) c58033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58033));
	wire w60033;

	wire w62033;
	repeater #(1, 1'b0, 0, 0) c62033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62033));
	wire w64033;

	wire w66033;
	repeater #(1, 1'b0, 0, 0) c66033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66033));
	wire w68033;

	wire w70033;
	repeater #(1, 1'b1, 0, 0) c70033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70033));
	wire w72033;

	wire w74033;
	repeater #(1, 1'b0, 0, 0) c74033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74033));
	wire w76033;

	wire w78033;
	repeater #(1, 1'b0, 0, 0) c78033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78033));
	wire w80033;

	wire w82033;
	repeater #(1, 1'b0, 0, 0) c82033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82033));
	wire w64037;
	torch #(1'b1) c64037 (.i_clk(tick), .i_in(), .o_out(w64037));
	wire w68037;
	torch #(1'b1) c68037 (.i_clk(tick), .i_in(), .o_out(w68037));
	wire w72037;
	torch #(1'b1) c72037 (.i_clk(tick), .i_in(), .o_out(w72037));
	wire w76037;
	torch #(1'b1) c76037 (.i_clk(tick), .i_in(), .o_out(w76037));
	wire w57046;
	torch #(1'b1) c57046 (.i_clk(tick), .i_in(), .o_out(w57046));
	wire w61046;
	torch #(1'b1) c61046 (.i_clk(tick), .i_in(), .o_out(w61046));
	wire w65046;
	torch #(1'b1) c65046 (.i_clk(tick), .i_in(), .o_out(w65046));
	wire w69046;
	torch #(1'b0) c69046 (.i_clk(tick), .i_in(), .o_out(w69046));
	wire w73046;
	torch #(1'b1) c73046 (.i_clk(tick), .i_in(), .o_out(w73046));
	wire w77046;
	torch #(1'b1) c77046 (.i_clk(tick), .i_in(), .o_out(w77046));
	wire w81046;
	torch #(1'b1) c81046 (.i_clk(tick), .i_in(), .o_out(w81046));
	wire w58047;
	repeater #(1, 1'b0, 0, 0) c58047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58047));
	wire w62047;
	repeater #(1, 1'b0, 0, 0) c62047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62047));
	wire w66047;
	repeater #(1, 1'b0, 0, 0) c66047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66047));
	wire w70047;
	repeater #(1, 1'b1, 0, 0) c70047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70047));
	wire w74047;
	repeater #(1, 1'b0, 0, 0) c74047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74047));
	wire w78047;
	repeater #(1, 1'b0, 0, 0) c78047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78047));
	wire w82047;
	repeater #(1, 1'b0, 0, 0) c82047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82047));
	wire w56049;

	wire w58049;
	repeater #(1, 1'b0, 0, 0) c58049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58049));
	wire w60049;

	wire w62049;
	repeater #(1, 1'b0, 0, 0) c62049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62049));
	wire w64049;

	wire w66049;
	repeater #(1, 1'b0, 0, 0) c66049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66049));
	wire w68049;

	wire w70049;
	repeater #(1, 1'b1, 0, 0) c70049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70049));
	wire w72049;

	wire w74049;
	repeater #(1, 1'b0, 0, 0) c74049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74049));
	wire w76049;

	wire w78049;
	repeater #(1, 1'b0, 0, 0) c78049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78049));
	wire w80049;

	wire w82049;
	repeater #(1, 1'b0, 0, 0) c82049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82049));
	wire w57055;
	torch #(1'b1) c57055 (.i_clk(tick), .i_in(), .o_out(w57055));
	wire w61055;
	torch #(1'b1) c61055 (.i_clk(tick), .i_in(), .o_out(w61055));
	wire w65055;
	torch #(1'b1) c65055 (.i_clk(tick), .i_in(), .o_out(w65055));
	wire w69055;
	torch #(1'b0) c69055 (.i_clk(tick), .i_in(), .o_out(w69055));
	wire w73055;
	torch #(1'b1) c73055 (.i_clk(tick), .i_in(), .o_out(w73055));
	wire w77055;
	torch #(1'b1) c77055 (.i_clk(tick), .i_in(), .o_out(w77055));
	wire w81055;
	torch #(1'b1) c81055 (.i_clk(tick), .i_in(), .o_out(w81055));
	wire w58067;
	repeater #(1, 1'b0, 0, 0) c58067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58067));
	wire w62067;
	repeater #(1, 1'b0, 0, 0) c62067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62067));
	wire w66067;
	repeater #(1, 1'b0, 0, 0) c66067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66067));
	wire w70067;
	repeater #(1, 1'b1, 0, 0) c70067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70067));
	wire w74067;
	repeater #(1, 1'b0, 0, 0) c74067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74067));
	wire w78067;
	repeater #(1, 1'b0, 0, 0) c78067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78067));
	wire w82067;
	repeater #(1, 1'b0, 0, 0) c82067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82067));
	wire w57068;
	repeater #(1, 1'b0, 0, 0) c57068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57068));
	wire w61068;
	repeater #(1, 1'b1, 0, 0) c61068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61068));
	wire w65068;
	repeater #(1, 1'b1, 0, 0) c65068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65068));
	wire w69068;
	repeater #(1, 1'b1, 0, 0) c69068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69068));
	wire w73068;
	repeater #(1, 1'b1, 0, 0) c73068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73068));
	wire w77068;
	repeater #(1, 1'b1, 0, 0) c77068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77068));
	wire w81068;
	repeater #(1, 1'b1, 0, 0) c81068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81068));
	wire w83074;
	repeater #(1, 1'b0, 0, 0) c83074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83074));
	wire w59077;
	repeater #(3, 1'b0, 0, 0) c59077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59077));
	wire w63077;
	repeater #(3, 1'b0, 0, 0) c63077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63077));
	wire w67077;
	repeater #(3, 1'b0, 0, 0) c67077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67077));
	wire w71077;
	repeater #(3, 1'b0, 0, 0) c71077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71077));
	wire w75077;
	repeater #(3, 1'b0, 0, 0) c75077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75077));
	wire w79077;
	repeater #(3, 1'b0, 0, 0) c79077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79077));
	wire w83077;
	repeater #(3, 1'b0, 0, 0) c83077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83077));
	wire w570102;
	torch #(1'b1) c570102 (.i_clk(tick), .i_in(), .o_out(w570102));
	wire w610102;
	torch #(1'b1) c610102 (.i_clk(tick), .i_in(), .o_out(w610102));
	wire w650102;
	torch #(1'b1) c650102 (.i_clk(tick), .i_in(), .o_out(w650102));
	wire w690102;
	torch #(1'b0) c690102 (.i_clk(tick), .i_in(), .o_out(w690102));
	wire w730102;
	torch #(1'b1) c730102 (.i_clk(tick), .i_in(), .o_out(w730102));
	wire w770102;
	torch #(1'b1) c770102 (.i_clk(tick), .i_in(), .o_out(w770102));
	wire w810102;
	torch #(1'b1) c810102 (.i_clk(tick), .i_in(), .o_out(w810102));
	wire w1730106;

	wire w2070106;

	wire w330107;

	wire w670107;

	wire w1720107;
	repeater #(1, 1'b1, 0, 0) c1720107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1720107));
	wire w2060107;
	repeater #(1, 1'b1, 0, 0) c2060107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060107));
	wire w320108;
	repeater #(1, 1'b1, 0, 0) c320108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320108));
	wire w660108;
	repeater #(1, 1'b1, 0, 0) c660108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660108));
	wire w1710108;

	wire w2050108;

	wire w310109;

	wire w650109;

	wire w1700109;
	repeater #(1, 1'b1, 0, 0) c1700109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1700109));
	wire w2040109;
	repeater #(1, 1'b1, 0, 0) c2040109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040109));
	wire w300110;
	repeater #(1, 1'b1, 0, 0) c300110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300110));
	wire w640110;
	repeater #(1, 1'b1, 0, 0) c640110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640110));
	wire w1690110;

	wire w2030110;

	wire w290111;

	wire w630111;

	wire w1680111;
	repeater #(1, 1'b1, 0, 0) c1680111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1680111));
	wire w2020111;
	repeater #(1, 1'b1, 0, 0) c2020111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020111));
	wire w280112;
	repeater #(1, 1'b1, 0, 0) c280112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280112));
	wire w620112;
	repeater #(1, 1'b1, 0, 0) c620112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620112));
	wire w1670112;

	wire w2010112;

	wire w270113;

	wire w610113;

	wire w1660113;
	repeater #(1, 1'b1, 0, 0) c1660113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1660113));
	wire w2000113;
	repeater #(1, 1'b1, 0, 0) c2000113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2000113));
	wire w260114;
	repeater #(1, 1'b1, 0, 0) c260114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260114));
	wire w600114;
	repeater #(1, 1'b1, 0, 0) c600114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600114));
	wire w1650114;

	wire w1990114;

	wire w250115;

	wire w590115;

	wire w1640115;
	repeater #(1, 1'b1, 0, 0) c1640115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640115));
	wire w1980115;
	repeater #(1, 1'b1, 0, 0) c1980115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980115));
	wire w240116;
	repeater #(1, 1'b1, 0, 0) c240116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240116));
	wire w580116;
	repeater #(1, 1'b1, 0, 0) c580116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580116));
	wire w1630116;

	wire w1970116;

	wire w230117;

	wire w570117;

	wire w1620117;
	repeater #(1, 1'b1, 0, 0) c1620117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620117));
	wire w1960117;
	repeater #(1, 1'b1, 0, 0) c1960117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1960117));
	wire w220118;
	repeater #(1, 1'b1, 0, 0) c220118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220118));
	wire w560118;
	repeater #(1, 1'b1, 0, 0) c560118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560118));
	wire w1610118;

	wire w1950118;

	wire w210119;

	wire w550119;

	wire w1600119;
	repeater #(1, 1'b1, 0, 0) c1600119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1600119));
	wire w1940119;
	repeater #(1, 1'b1, 0, 0) c1940119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1940119));
	wire w200120;
	repeater #(1, 1'b1, 0, 0) c200120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200120));
	wire w540120;
	repeater #(1, 1'b1, 0, 0) c540120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540120));
	wire w1590120;

	wire w1930120;

	wire w190121;

	wire w530121;

	wire w1580121;
	repeater #(1, 1'b0, 0, 0) c1580121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580121));
	wire w1920121;
	repeater #(1, 1'b0, 0, 0) c1920121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1920121));
	wire w180122;
	repeater #(1, 1'b0, 0, 0) c180122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180122));
	wire w520122;
	repeater #(1, 1'b0, 0, 0) c520122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520122));
	wire w1570122;

	wire w1910122;

	wire w170123;

	wire w510123;

	wire w1560123;
	repeater #(1, 1'b1, 0, 0) c1560123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560123));
	wire w1900123;
	repeater #(1, 1'b1, 0, 0) c1900123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1900123));
	wire w160124;
	repeater #(1, 1'b1, 0, 0) c160124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160124));
	wire w500124;
	repeater #(1, 1'b1, 0, 0) c500124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500124));
	wire w1550124;

	wire w1890124;

	wire w150125;

	wire w490125;

	wire w1540125;
	repeater #(1, 1'b1, 0, 0) c1540125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540125));
	wire w1880125;
	repeater #(1, 1'b1, 0, 0) c1880125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1880125));
	wire w140126;
	repeater #(1, 1'b1, 0, 0) c140126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140126));
	wire w480126;
	repeater #(1, 1'b1, 0, 0) c480126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480126));
	wire w1530126;

	wire w1870126;

	wire w130127;

	wire w470127;

	wire w1520127;
	repeater #(1, 1'b1, 0, 0) c1520127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520127));
	wire w1860127;
	repeater #(1, 1'b1, 0, 0) c1860127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860127));
	wire w120128;
	repeater #(1, 1'b1, 0, 0) c120128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120128));
	wire w460128;
	repeater #(1, 1'b1, 0, 0) c460128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460128));
	wire w1510128;

	wire w1850128;

	wire w110129;

	wire w450129;

	wire w1500129;
	repeater #(1, 1'b1, 0, 0) c1500129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500129));
	wire w1840129;
	repeater #(1, 1'b1, 0, 0) c1840129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1840129));
	wire w100130;
	repeater #(1, 1'b1, 0, 0) c100130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100130));
	wire w440130;
	repeater #(1, 1'b1, 0, 0) c440130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440130));
	wire w1490130;

	wire w1830130;

	wire w90131;

	wire w430131;

	wire w1480131;
	repeater #(1, 1'b1, 0, 0) c1480131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1480131));
	wire w1820131;
	repeater #(1, 1'b1, 0, 0) c1820131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820131));
	wire w80132;
	repeater #(1, 1'b1, 0, 0) c80132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80132));
	wire w420132;
	repeater #(1, 1'b1, 0, 0) c420132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420132));
	wire w1470132;

	wire w1810132;

	wire w70133;

	wire w410133;

	wire w1460133;
	repeater #(1, 1'b1, 0, 0) c1460133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460133));
	wire w1800133;
	repeater #(1, 1'b1, 0, 0) c1800133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800133));
	wire w60134;
	repeater #(1, 1'b1, 0, 0) c60134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60134));
	wire w400134;
	repeater #(1, 1'b1, 0, 0) c400134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400134));
	wire w1440138;
	repeater #(2, 1'b1, 0, 0) c1440138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1440138));
	wire w1780138;
	repeater #(2, 1'b1, 0, 0) c1780138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1780138));
	wire w560140;
	repeater #(1, 1'b1, 0, 0) c560140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560140));
	wire w600140;
	repeater #(1, 1'b1, 0, 0) c600140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600140));
	wire w640140;
	repeater #(1, 1'b1, 0, 0) c640140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640140));
	wire w680140;
	repeater #(1, 1'b0, 0, 0) c680140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w680140));
	wire w720140;
	repeater #(1, 1'b1, 0, 0) c720140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w720140));
	wire w760140;
	repeater #(1, 1'b1, 0, 0) c760140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w760140));
	wire w800140;
	repeater #(1, 1'b1, 0, 0) c800140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800140));
	wire w1300140;
	repeater #(1, 1'b1, 0, 0) c1300140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1300140));
	wire w1360140;
	torch #(1'b1) c1360140 (.i_clk(tick), .i_in(), .o_out(w1360140));
	wire w1460140;
	repeater #(1, 1'b1, 0, 0) c1460140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460140));
	wire w1520140;
	torch #(1'b0) c1520140 (.i_clk(tick), .i_in(), .o_out(w1520140));
	wire w1640140;
	repeater #(1, 1'b1, 0, 0) c1640140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640140));
	wire w1700140;
	torch #(1'b1) c1700140 (.i_clk(tick), .i_in(), .o_out(w1700140));
	wire w1800140;
	repeater #(1, 1'b1, 0, 0) c1800140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800140));
	wire w1860140;
	torch #(1'b0) c1860140 (.i_clk(tick), .i_in(), .o_out(w1860140));
	wire w560141;
	repeater #(1, 1'b1, 0, 0) c560141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560141));
	wire w580141;
	repeater #(1, 1'b0, 0, 0) c580141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580141));
	wire w600141;
	repeater #(1, 1'b1, 0, 0) c600141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600141));
	wire w620141;
	repeater #(1, 1'b0, 0, 0) c620141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620141));
	wire w640141;
	repeater #(1, 1'b1, 0, 0) c640141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640141));
	wire w660141;
	repeater #(1, 1'b0, 0, 0) c660141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660141));
	wire w680141;
	repeater #(1, 1'b0, 0, 0) c680141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w680141));
	wire w700141;
	repeater #(1, 1'b0, 0, 0) c700141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w700141));
	wire w720141;
	repeater #(1, 1'b1, 0, 0) c720141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w720141));
	wire w740141;
	repeater #(1, 1'b0, 0, 0) c740141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w740141));
	wire w760141;
	repeater #(1, 1'b1, 0, 0) c760141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w760141));
	wire w780141;
	repeater #(1, 1'b0, 0, 0) c780141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w780141));
	wire w800141;
	repeater #(1, 1'b1, 0, 0) c800141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800141));
	wire w820141;
	repeater #(1, 1'b0, 0, 0) c820141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w820141));
	wire w570142;
	torch #(1'b0) c570142 (.i_clk(tick), .i_in(), .o_out(w570142));
	wire w610142;
	torch #(1'b0) c610142 (.i_clk(tick), .i_in(), .o_out(w610142));
	wire w650142;
	torch #(1'b0) c650142 (.i_clk(tick), .i_in(), .o_out(w650142));
	wire w690142;
	torch #(1'b0) c690142 (.i_clk(tick), .i_in(), .o_out(w690142));
	wire w730142;
	torch #(1'b0) c730142 (.i_clk(tick), .i_in(), .o_out(w730142));
	wire w770142;
	torch #(1'b0) c770142 (.i_clk(tick), .i_in(), .o_out(w770142));
	wire w810142;
	torch #(1'b0) c810142 (.i_clk(tick), .i_in(), .o_out(w810142));
	wire w1370143;
	repeater #(1, 1'b1, 0, 0) c1370143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370143));
	wire w1530143;
	repeater #(1, 1'b0, 0, 0) c1530143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1530143));
	wire w1710143;
	repeater #(1, 1'b1, 0, 0) c1710143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710143));
	wire w1870143;
	repeater #(1, 1'b1, 0, 0) c1870143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870143));
	wire w1300144;
	repeater #(1, 1'b1, 0, 0) c1300144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1300144));
	wire w1460144;
	repeater #(1, 1'b1, 0, 0) c1460144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460144));
	wire w1640144;
	repeater #(1, 1'b1, 0, 0) c1640144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640144));
	wire w1800144;
	repeater #(1, 1'b1, 0, 0) c1800144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800144));
	wire w2050144;
	repeater #(1, 1'b0, 0, 0) c2050144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2050144));
	wire w10145;
	repeater #(1, 1'b0, 0, 0) c10145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10145));
	wire w50145;
	repeater #(1, 1'b0, 0, 0) c50145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50145));
	wire w90145;
	repeater #(1, 1'b0, 0, 0) c90145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90145));
	wire w290145;
	repeater #(1, 1'b1, 0, 0) c290145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290145));
	wire w330145;
	repeater #(1, 1'b1, 0, 0) c330145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330145));
	wire w370145;
	repeater #(1, 1'b1, 0, 0) c370145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370145));
	wire w410145;
	repeater #(1, 1'b1, 0, 0) c410145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w410145));
	wire w1350145;

	wire w1510145;

	wire w1690145;

	wire w1850145;

	wire w1430146;

	wire w1770146;

	wire w1290147;

	wire w1300147;

	wire w1400147;

	wire w1450147;

	wire w1460147;

	wire w1630147;

	wire w1640147;

	wire w1740147;

	wire w1790147;

	wire w1800147;

	wire w2030147;
	torch #(1'b0) c2030147 (.i_clk(tick), .i_in(), .o_out(w2030147));
	wire w2070147;
	torch #(1'b1) c2070147 (.i_clk(tick), .i_in(), .o_out(w2070147));
	wire w30148;
	torch #(1'b1) c30148 (.i_clk(tick), .i_in(), .o_out(w30148));
	wire w70148;
	torch #(1'b0) c70148 (.i_clk(tick), .i_in(), .o_out(w70148));
	wire w310148;
	torch #(1'b1) c310148 (.i_clk(tick), .i_in(), .o_out(w310148));
	wire w350148;
	torch #(1'b0) c350148 (.i_clk(tick), .i_in(), .o_out(w350148));
	wire w390148;
	torch #(1'b0) c390148 (.i_clk(tick), .i_in(), .o_out(w390148));
	wire w430148;
	torch #(1'b0) c430148 (.i_clk(tick), .i_in(), .o_out(w430148));
	wire w640149;
	torch #(1'b1) c640149 (.i_clk(tick), .i_in(), .o_out(w640149));
	wire w680149;
	torch #(1'b1) c680149 (.i_clk(tick), .i_in(), .o_out(w680149));
	wire w720149;
	torch #(1'b1) c720149 (.i_clk(tick), .i_in(), .o_out(w720149));
	wire w760149;
	torch #(1'b1) c760149 (.i_clk(tick), .i_in(), .o_out(w760149));
	wire w1380149;

	wire w1720149;

	wire w1280150;

	wire w1290150;

	wire w1440150;

	wire w1450150;

	wire w1620150;

	wire w1630150;

	wire w1780150;

	wire w1790150;

	wire w1300151;

	wire w1340151;

	wire w1380151;

	wire w1640151;

	wire w1680151;

	wire w1720151;

	wire w580152;

	wire w620152;

	wire w660152;

	wire w700152;

	wire w740152;

	wire w780152;

	wire w820152;

	wire w1540154;

	wire w1880154;

	wire w1270155;

	wire w1280155;

	wire w1310155;

	wire w1320155;

	wire w1350155;

	wire w1360155;

	wire w1390155;

	wire w1400155;

	wire w1430155;

	wire w1440155;

	wire w1470155;

	wire w1480155;

	wire w1510155;

	wire w1520155;

	wire w1610155;

	wire w1620155;

	wire w1650155;

	wire w1660155;

	wire w1690155;

	wire w1700155;

	wire w1730155;

	wire w1740155;

	wire w1770155;

	wire w1780155;

	wire w1810155;

	wire w1820155;

	wire w1850155;

	wire w1860155;

	wire w1250156;

	wire w1590156;

	wire w1400159;
	repeater #(1, 1'b1, 0, 0) c1400159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1400159));
	wire w1440159;
	repeater #(1, 1'b1, 0, 0) c1440159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1440159));
	wire w1480159;
	repeater #(1, 1'b1, 0, 0) c1480159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1480159));
	wire w1740159;
	repeater #(1, 1'b1, 0, 0) c1740159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1740159));
	wire w1780159;
	repeater #(1, 1'b1, 0, 0) c1780159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1780159));
	wire w1820159;
	repeater #(1, 1'b1, 0, 0) c1820159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820159));
	wire w1260162;

	wire w1300162;

	wire w1460162;

	wire w1500162;

	wire w1600162;

	wire w1640162;

	wire w1800162;

	wire w1840162;

	wire w580163;
	torch #(1'b0) c580163 (.i_clk(tick), .i_in(), .o_out(w580163));
	wire w620163;
	torch #(1'b0) c620163 (.i_clk(tick), .i_in(), .o_out(w620163));
	wire w660163;
	torch #(1'b0) c660163 (.i_clk(tick), .i_in(), .o_out(w660163));
	wire w700163;
	torch #(1'b1) c700163 (.i_clk(tick), .i_in(), .o_out(w700163));
	wire w740163;
	torch #(1'b0) c740163 (.i_clk(tick), .i_in(), .o_out(w740163));
	wire w780163;
	torch #(1'b0) c780163 (.i_clk(tick), .i_in(), .o_out(w780163));
	wire w820163;
	torch #(1'b0) c820163 (.i_clk(tick), .i_in(), .o_out(w820163));
	wire w1280163;
	repeater #(1, 1'b1, 0, 0) c1280163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1280163));
	wire w1440163;
	repeater #(1, 1'b1, 0, 0) c1440163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1440163));
	wire w1620163;
	repeater #(1, 1'b1, 0, 0) c1620163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620163));
	wire w1780163;
	repeater #(1, 1'b1, 0, 0) c1780163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1780163));
	wire w1220164;

	wire w1350164;
	repeater #(1, 1'b0, 0, 0) c1350164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350164));
	wire w1560164;

	wire w1690164;
	repeater #(1, 1'b1, 0, 0) c1690164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1690164));
	wire w640165;
	torch #(1'b1) c640165 (.i_clk(tick), .i_in(), .o_out(w640165));
	wire w680165;
	torch #(1'b1) c680165 (.i_clk(tick), .i_in(), .o_out(w680165));
	wire w720165;
	torch #(1'b1) c720165 (.i_clk(tick), .i_in(), .o_out(w720165));
	wire w760165;
	torch #(1'b1) c760165 (.i_clk(tick), .i_in(), .o_out(w760165));
	wire w1300165;

	wire w1460165;

	wire w1640165;

	wire w1800165;

	wire w1220166;

	wire w1380166;

	wire w1560166;

	wire w1720166;

	wire w1250167;

	wire w1330167;

	wire w1350167;

	wire w1360167;

	wire w1410167;

	wire w1490167;

	wire w1590167;

	wire w1670167;

	wire w1690167;

	wire w1700167;

	wire w1750167;

	wire w1830167;

	wire w580168;

	wire w620168;

	wire w660168;

	wire w700168;

	wire w740168;

	wire w780168;

	wire w820168;

	wire w1270169;

	wire w1280169;

	wire w1430169;

	wire w1440169;

	wire w1610169;

	wire w1620169;

	wire w1770169;

	wire w1780169;

	wire w100170;
	repeater #(1, 1'b0, 0, 0) c100170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100170));
	wire w280170;
	repeater #(1, 1'b1, 0, 0) c280170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280170));
	wire w1330171;

	wire w1350171;

	wire w1360171;

	wire w1490171;

	wire w1670171;

	wire w1690171;

	wire w1700171;

	wire w1830171;

	wire w180172;

	wire w170173;
	repeater #(1, 1'b0, 0, 0) c170173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170173));
	wire w1300173;
	torch #(1'b1) c1300173 (.i_clk(tick), .i_in(), .o_out(w1300173));
	wire w1310173;

	wire w1460173;
	torch #(1'b1) c1460173 (.i_clk(tick), .i_in(), .o_out(w1460173));
	wire w1470173;

	wire w1640173;
	torch #(1'b1) c1640173 (.i_clk(tick), .i_in(), .o_out(w1640173));
	wire w1650173;

	wire w1800173;
	torch #(1'b1) c1800173 (.i_clk(tick), .i_in(), .o_out(w1800173));
	wire w1810173;

	wire w1310174;

	wire w1330174;

	wire w1470174;

	wire w1490174;

	wire w1650174;

	wire w1670174;

	wire w1810174;

	wire w1830174;

	wire w210175;

	wire w180176;

	wire w1330176;

	wire w1340176;

	wire w1350176;

	wire w1490176;

	wire w1500176;

	wire w1510176;

	wire w1670176;

	wire w1680176;

	wire w1690176;

	wire w1830176;

	wire w1840176;

	wire w1850176;

	wire w2070176;

	wire w30177;
	repeater #(1, 1'b0, 0, 0) c30177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30177));
	wire w170177;

	wire w190177;
	repeater #(2, 1'b0, 0, 0) c190177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190177));
	wire w220177;
	repeater #(2, 1'b0, 0, 0) c220177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220177));
	wire w350177;
	repeater #(1, 1'b0, 0, 0) c350177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w350177));
	wire w390177;

	wire w1280177;

	wire w1290177;

	wire w1350177;

	wire w1440177;

	wire w1450177;

	wire w1510177;

	wire w1620177;

	wire w1630177;

	wire w1690177;

	wire w1780177;

	wire w1790177;

	wire w1850177;

	wire w00178;

	wire w60178;
	repeater #(2, 1'b0, 0, 0) c60178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60178));
	wire w90178;
	repeater #(2, 1'b1, 0, 0) c90178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90178));
	wire w110178;

	wire w270178;

	wire w290178;
	repeater #(2, 1'b0, 0, 0) c290178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290178));
	wire w320178;
	repeater #(2, 1'b0, 0, 0) c320178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320178));
	wire w380178;

	wire w1010;

	wire w2810;

	wire w5810;
	torch #(1'b0) c5810 (.i_clk(tick), .i_in(), .o_out(w5810));
	wire w6210;
	torch #(1'b0) c6210 (.i_clk(tick), .i_in(), .o_out(w6210));
	wire w6610;
	torch #(1'b0) c6610 (.i_clk(tick), .i_in(), .o_out(w6610));
	wire w7010;
	torch #(1'b1) c7010 (.i_clk(tick), .i_in(), .o_out(w7010));
	wire w7410;
	torch #(1'b0) c7410 (.i_clk(tick), .i_in(), .o_out(w7410));
	wire w7810;
	torch #(1'b0) c7810 (.i_clk(tick), .i_in(), .o_out(w7810));
	wire w8210;
	torch #(1'b0) c8210 (.i_clk(tick), .i_in(), .o_out(w8210));
	wire w13310;
	repeater #(1, 1'b0, 0, 0) c13310 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13310));
	wire w13510;
	torch #(1'b0) c13510 (.i_clk(tick), .i_in(), .o_out(w13510));
	wire w14110;
	torch #(1'b1) c14110 (.i_clk(tick), .i_in(), .o_out(w14110));
	wire w14910;
	repeater #(1, 1'b0, 0, 0) c14910 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14910));
	wire w15110;
	torch #(1'b0) c15110 (.i_clk(tick), .i_in(), .o_out(w15110));
	wire w16710;
	repeater #(1, 1'b0, 0, 0) c16710 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16710));
	wire w16910;
	torch #(1'b0) c16910 (.i_clk(tick), .i_in(), .o_out(w16910));
	wire w17510;
	torch #(1'b1) c17510 (.i_clk(tick), .i_in(), .o_out(w17510));
	wire w18310;
	repeater #(1, 1'b0, 0, 0) c18310 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18310));
	wire w18510;
	torch #(1'b0) c18510 (.i_clk(tick), .i_in(), .o_out(w18510));
	wire w711;

	wire w3111;

	wire w6412;
	torch #(1'b1) c6412 (.i_clk(tick), .i_in(), .o_out(w6412));
	wire w6812;
	torch #(1'b1) c6812 (.i_clk(tick), .i_in(), .o_out(w6812));
	wire w7212;
	torch #(1'b1) c7212 (.i_clk(tick), .i_in(), .o_out(w7212));
	wire w7612;
	torch #(1'b1) c7612 (.i_clk(tick), .i_in(), .o_out(w7612));
	wire w13712;
	repeater #(1, 1'b1, 0, 0) c13712 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13712));
	wire w15312;
	repeater #(1, 1'b1, 0, 0) c15312 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15312));
	wire w17112;
	repeater #(1, 1'b1, 0, 0) c17112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17112));
	wire w18712;
	repeater #(1, 1'b1, 0, 0) c18712 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18712));
	wire w2513;
	assign outputs[38] = ();
	wire w13414;
	torch #(1'b1) c13414 (.i_clk(tick), .i_in(), .o_out(w13414));
	wire w15014;
	torch #(1'b1) c15014 (.i_clk(tick), .i_in(), .o_out(w15014));
	wire w16814;
	torch #(1'b1) c16814 (.i_clk(tick), .i_in(), .o_out(w16814));
	wire w18414;
	torch #(1'b1) c18414 (.i_clk(tick), .i_in(), .o_out(w18414));
	wire w5815;

	wire w6215;

	wire w6615;

	wire w7015;

	wire w7415;

	wire w7815;

	wire w8215;

	wire w14216;
	torch #(1'b1) c14216 (.i_clk(tick), .i_in(), .o_out(w14216));
	wire w17616;
	torch #(1'b1) c17616 (.i_clk(tick), .i_in(), .o_out(w17616));
	wire w13317;
	repeater #(2, 1'b0, 0, 0) c13317 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13317));
	wire w14917;
	repeater #(1, 1'b0, 0, 0) c14917 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14917));
	wire w16717;
	repeater #(2, 1'b0, 0, 0) c16717 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16717));
	wire w18317;
	repeater #(1, 1'b0, 0, 0) c18317 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18317));
	wire w14318;
	repeater #(1, 1'b0, 0, 0) c14318 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14318));
	wire w17718;
	repeater #(1, 1'b0, 0, 0) c17718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17718));
	wire w137110;
	repeater #(1, 1'b0, 0, 0) c137110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137110));
	wire w171110;
	repeater #(1, 1'b0, 0, 0) c171110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171110));
	wire w139111;
	repeater #(1, 1'b0, 0, 0) c139111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139111));
	wire w173111;
	repeater #(1, 1'b0, 0, 0) c173111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173111));
	wire w58116;
	torch #(1'b0) c58116 (.i_clk(tick), .i_in(), .o_out(w58116));
	wire w62116;
	torch #(1'b0) c62116 (.i_clk(tick), .i_in(), .o_out(w62116));
	wire w66116;
	torch #(1'b0) c66116 (.i_clk(tick), .i_in(), .o_out(w66116));
	wire w70116;
	torch #(1'b1) c70116 (.i_clk(tick), .i_in(), .o_out(w70116));
	wire w74116;
	torch #(1'b0) c74116 (.i_clk(tick), .i_in(), .o_out(w74116));
	wire w78116;
	torch #(1'b0) c78116 (.i_clk(tick), .i_in(), .o_out(w78116));
	wire w82116;
	torch #(1'b0) c82116 (.i_clk(tick), .i_in(), .o_out(w82116));
	wire w64118;
	torch #(1'b1) c64118 (.i_clk(tick), .i_in(), .o_out(w64118));
	wire w68118;
	torch #(1'b1) c68118 (.i_clk(tick), .i_in(), .o_out(w68118));
	wire w72118;
	torch #(1'b1) c72118 (.i_clk(tick), .i_in(), .o_out(w72118));
	wire w76118;
	torch #(1'b1) c76118 (.i_clk(tick), .i_in(), .o_out(w76118));
	wire w58121;

	wire w62121;

	wire w66121;

	wire w70121;

	wire w74121;

	wire w78121;

	wire w82121;

	wire w12125;

	wire w30125;

	wire w58132;
	torch #(1'b0) c58132 (.i_clk(tick), .i_in(), .o_out(w58132));
	wire w62132;
	torch #(1'b0) c62132 (.i_clk(tick), .i_in(), .o_out(w62132));
	wire w66132;
	torch #(1'b0) c66132 (.i_clk(tick), .i_in(), .o_out(w66132));
	wire w70132;
	torch #(1'b1) c70132 (.i_clk(tick), .i_in(), .o_out(w70132));
	wire w74132;
	torch #(1'b0) c74132 (.i_clk(tick), .i_in(), .o_out(w74132));
	wire w78132;
	torch #(1'b0) c78132 (.i_clk(tick), .i_in(), .o_out(w78132));
	wire w82132;
	torch #(1'b0) c82132 (.i_clk(tick), .i_in(), .o_out(w82132));
	wire w64134;
	torch #(1'b1) c64134 (.i_clk(tick), .i_in(), .o_out(w64134));
	wire w68134;
	torch #(1'b1) c68134 (.i_clk(tick), .i_in(), .o_out(w68134));
	wire w72134;
	torch #(1'b1) c72134 (.i_clk(tick), .i_in(), .o_out(w72134));
	wire w76134;
	torch #(1'b1) c76134 (.i_clk(tick), .i_in(), .o_out(w76134));
	wire w58137;

	wire w62137;

	wire w66137;

	wire w70137;

	wire w74137;

	wire w78137;

	wire w82137;

	wire w58148;
	torch #(1'b0) c58148 (.i_clk(tick), .i_in(), .o_out(w58148));
	wire w62148;
	torch #(1'b0) c62148 (.i_clk(tick), .i_in(), .o_out(w62148));
	wire w66148;
	torch #(1'b0) c66148 (.i_clk(tick), .i_in(), .o_out(w66148));
	wire w70148;
	torch #(1'b1) c70148 (.i_clk(tick), .i_in(), .o_out(w70148));
	wire w74148;
	torch #(1'b0) c74148 (.i_clk(tick), .i_in(), .o_out(w74148));
	wire w78148;
	torch #(1'b0) c78148 (.i_clk(tick), .i_in(), .o_out(w78148));
	wire w82148;
	torch #(1'b0) c82148 (.i_clk(tick), .i_in(), .o_out(w82148));
	wire w56151;
	assign outputs[39] = ();
	wire w58151;
	assign outputs[40] = ();
	wire w60151;
	assign outputs[41] = ();
	wire w62151;
	assign outputs[42] = ();
	wire w64151;
	assign outputs[43] = ();
	wire w66151;
	assign outputs[44] = ();
	wire w68151;
	assign outputs[45] = ();
	wire w70151;
	assign outputs[46] = ();
	wire w72151;
	assign outputs[47] = ();
	wire w74151;
	assign outputs[48] = ();
	wire w76151;
	assign outputs[49] = ();
	wire w78151;
	assign outputs[50] = ();
	wire w80151;
	assign outputs[51] = ();
	wire w82151;
	assign outputs[52] = ();
	wire w56152;
	repeater #(1, 1'b0, 0, 0) c56152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56152));
	wire w58152;
	repeater #(1, 1'b0, 0, 0) c58152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58152));
	wire w60152;
	repeater #(1, 1'b0, 0, 0) c60152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60152));
	wire w62152;
	repeater #(1, 1'b0, 0, 0) c62152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62152));
	wire w64152;
	repeater #(1, 1'b0, 0, 0) c64152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64152));
	wire w66152;
	repeater #(1, 1'b0, 0, 0) c66152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66152));
	wire w68152;
	repeater #(1, 1'b0, 0, 0) c68152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68152));
	wire w70152;
	repeater #(1, 1'b1, 0, 0) c70152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70152));
	wire w72152;
	repeater #(1, 1'b0, 0, 0) c72152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72152));
	wire w74152;
	repeater #(1, 1'b0, 0, 0) c74152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74152));
	wire w76152;
	repeater #(1, 1'b0, 0, 0) c76152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76152));
	wire w78152;
	repeater #(1, 1'b0, 0, 0) c78152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78152));
	wire w80152;
	repeater #(1, 1'b0, 0, 0) c80152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80152));
	wire w82152;
	repeater #(1, 1'b0, 0, 0) c82152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82152));
	wire w57159;
	repeater #(2, 1'b1, 0, 0) c57159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57159));
	wire w61159;
	repeater #(2, 1'b1, 0, 0) c61159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61159));
	wire w65159;
	repeater #(2, 1'b1, 0, 0) c65159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65159));
	wire w69159;
	repeater #(2, 1'b0, 0, 0) c69159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69159));
	wire w73159;
	repeater #(2, 1'b1, 0, 0) c73159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73159));
	wire w77159;
	repeater #(2, 1'b1, 0, 0) c77159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77159));
	wire w81159;
	repeater #(2, 1'b1, 0, 0) c81159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81159));
	wire w55164;
	repeater #(1, 1'b1, 0, 0) c55164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55164));
	wire w59164;
	repeater #(1, 1'b1, 0, 0) c59164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59164));
	wire w63164;
	repeater #(1, 1'b1, 0, 0) c63164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63164));
	wire w67164;
	repeater #(1, 1'b0, 0, 0) c67164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67164));
	wire w71164;
	repeater #(1, 1'b1, 0, 0) c71164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71164));
	wire w75164;
	repeater #(1, 1'b1, 0, 0) c75164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75164));
	wire w79164;
	repeater #(1, 1'b1, 0, 0) c79164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79164));
	wire w57165;

	wire w61165;

	wire w65165;

	wire w69165;

	wire w73165;

	wire w77165;

	wire w81165;

	wire w56166;

	wire w60166;

	wire w64166;

	wire w68166;

	wire w72166;

	wire w76166;

	wire w80166;

	wire w57167;
	torch #(1'b1) c57167 (.i_clk(tick), .i_in(), .o_out(w57167));
	wire w61167;
	torch #(1'b1) c61167 (.i_clk(tick), .i_in(), .o_out(w61167));
	wire w65167;
	torch #(1'b1) c65167 (.i_clk(tick), .i_in(), .o_out(w65167));
	wire w69167;
	torch #(1'b1) c69167 (.i_clk(tick), .i_in(), .o_out(w69167));
	wire w73167;
	torch #(1'b1) c73167 (.i_clk(tick), .i_in(), .o_out(w73167));
	wire w77167;
	torch #(1'b1) c77167 (.i_clk(tick), .i_in(), .o_out(w77167));
	wire w81167;
	torch #(1'b1) c81167 (.i_clk(tick), .i_in(), .o_out(w81167));
	wire w55168;
	repeater #(1, 1'b1, 0, 0) c55168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55168));
	wire w59168;
	repeater #(1, 1'b1, 0, 0) c59168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59168));
	wire w63168;
	repeater #(1, 1'b1, 0, 0) c63168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63168));
	wire w67168;
	repeater #(1, 1'b1, 0, 0) c67168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67168));
	wire w71168;
	repeater #(1, 1'b1, 0, 0) c71168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71168));
	wire w75168;
	repeater #(1, 1'b1, 0, 0) c75168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75168));
	wire w79168;
	repeater #(1, 1'b1, 0, 0) c79168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79168));
	wire w72172;
	torch #(1'b0) c72172 (.i_clk(tick), .i_in(), .o_out(w72172));
	wire w57180;
	assign w57180 = inputs[13];
	wire w61180;
	assign w61180 = inputs[14];
	wire w65180;
	assign w65180 = inputs[15];
	wire w69180;
	assign w69180 = inputs[16];
	wire w73180;
	assign w73180 = inputs[17];
	wire w77180;
	assign w77180 = inputs[18];
	wire w81180;
	assign w81180 = inputs[19];
	wire w821126;

	wire w801128;

	wire w781130;

	wire w761132;

	wire w741134;

	wire w12402;
	repeater #(2, 1'b0, 0, 0) c12402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12402));
	wire w15802;
	repeater #(2, 1'b0, 0, 0) c15802 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15802));
	wire w4104;
	torch #(1'b1) c4104 (.i_clk(tick), .i_in(), .o_out(w4104));
	wire w4504;
	torch #(1'b1) c4504 (.i_clk(tick), .i_in(), .o_out(w4504));
	wire w4904;
	torch #(1'b1) c4904 (.i_clk(tick), .i_in(), .o_out(w4904));
	wire w5304;
	torch #(1'b1) c5304 (.i_clk(tick), .i_in(), .o_out(w5304));
	wire w5704;
	torch #(1'b1) c5704 (.i_clk(tick), .i_in(), .o_out(w5704));
	wire w6104;
	torch #(1'b1) c6104 (.i_clk(tick), .i_in(), .o_out(w6104));
	wire w6504;
	torch #(1'b1) c6504 (.i_clk(tick), .i_in(), .o_out(w6504));
	wire w11604;
	torch #(1'b1) c11604 (.i_clk(tick), .i_in(), .o_out(w11604));
	wire w12604;
	repeater #(1, 1'b0, 0, 0) c12604 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12604));
	wire w13204;
	torch #(1'b1) c13204 (.i_clk(tick), .i_in(), .o_out(w13204));
	wire w15004;
	torch #(1'b1) c15004 (.i_clk(tick), .i_in(), .o_out(w15004));
	wire w16004;
	repeater #(1, 1'b1, 0, 0) c16004 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16004));
	wire w16604;
	torch #(1'b1) c16604 (.i_clk(tick), .i_in(), .o_out(w16604));
	wire w4207;
	repeater #(2, 1'b0, 0, 0) c4207 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4207));
	wire w4607;
	repeater #(2, 1'b0, 0, 0) c4607 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4607));
	wire w5007;
	repeater #(2, 1'b0, 0, 0) c5007 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5007));
	wire w5407;
	repeater #(2, 1'b0, 0, 0) c5407 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5407));
	wire w5807;
	repeater #(1, 1'b0, 0, 0) c5807 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5807));
	wire w6207;
	repeater #(1, 1'b0, 0, 0) c6207 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6207));
	wire w6607;
	repeater #(1, 1'b0, 0, 0) c6607 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6607));
	wire w11707;
	repeater #(1, 1'b1, 0, 0) c11707 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11707));
	wire w13307;
	repeater #(1, 1'b1, 0, 0) c13307 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13307));
	wire w15107;
	repeater #(1, 1'b1, 0, 0) c15107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15107));
	wire w16707;
	repeater #(1, 1'b1, 0, 0) c16707 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16707));
	wire w5508;
	repeater #(1, 1'b0, 0, 0) c5508 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5508));
	wire w6708;
	repeater #(2, 1'b0, 0, 0) c6708 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6708));
	wire w12608;
	repeater #(1, 1'b0, 0, 0) c12608 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12608));
	wire w13908;

	wire w16008;
	repeater #(1, 1'b1, 0, 0) c16008 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16008));
	wire w17308;

	wire w11509;

	wire w13109;

	wire w14909;

	wire w16509;

	wire w123010;

	wire w139010;

	wire w157010;

	wire w173010;

	wire w120011;

	wire w125011;

	wire w126011;

	wire w136011;

	wire w154011;

	wire w159011;

	wire w160011;

	wire w170011;

	wire w44013;
	repeater #(1, 1'b0, 0, 0) c44013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44013));
	wire w64013;
	repeater #(1, 1'b0, 0, 0) c64013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64013));
	wire w118013;

	wire w134013;

	wire w152013;

	wire w168013;

	wire w124014;

	wire w125014;

	wire w158014;

	wire w159014;

	wire w110015;

	wire w144015;

	wire w189015;
	repeater #(1, 1'b1, 0, 0) c189015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189015));
	wire w191015;
	repeater #(2, 1'b1, 0, 0) c191015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191015));
	wire w193015;
	repeater #(2, 1'b0, 0, 0) c193015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193015));
	wire w197015;
	repeater #(2, 1'b0, 0, 0) c197015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197015));
	wire w199015;
	repeater #(2, 1'b1, 0, 0) c199015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199015));
	wire w201015;
	repeater #(1, 1'b1, 0, 0) c201015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201015));
	wire w13016;
	repeater #(1, 1'b1, 0, 0) c13016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13016));
	wire w15016;
	repeater #(2, 1'b0, 0, 0) c15016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15016));
	wire w17016;
	repeater #(2, 1'b1, 0, 0) c17016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17016));
	wire w21016;
	repeater #(2, 1'b1, 0, 0) c21016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21016));
	wire w23016;
	repeater #(2, 1'b1, 0, 0) c23016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23016));
	wire w25016;
	repeater #(1, 1'b1, 0, 0) c25016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25016));
	wire w186016;
	repeater #(1, 1'b1, 0, 0) c186016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186016));
	wire w28017;
	repeater #(1, 1'b1, 0, 0) c28017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28017));
	wire w111017;
	repeater #(1, 1'b1, 0, 0) c111017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111017));
	wire w115017;
	repeater #(1, 1'b1, 0, 0) c115017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115017));
	wire w119017;
	repeater #(1, 1'b1, 0, 0) c119017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119017));
	wire w123017;
	repeater #(1, 1'b0, 0, 0) c123017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123017));
	wire w127017;
	repeater #(1, 1'b1, 0, 0) c127017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127017));
	wire w131017;
	repeater #(1, 1'b1, 0, 0) c131017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131017));
	wire w135017;
	repeater #(1, 1'b1, 0, 0) c135017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135017));
	wire w145017;
	repeater #(1, 1'b1, 0, 0) c145017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145017));
	wire w149017;
	repeater #(1, 1'b1, 0, 0) c149017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149017));
	wire w153017;
	repeater #(1, 1'b1, 0, 0) c153017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153017));
	wire w157017;
	repeater #(1, 1'b1, 0, 0) c157017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157017));
	wire w161017;
	repeater #(1, 1'b1, 0, 0) c161017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161017));
	wire w165017;
	repeater #(1, 1'b1, 0, 0) c165017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165017));
	wire w169017;
	repeater #(1, 1'b1, 0, 0) c169017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169017));
	wire w196017;

	wire w18018;

	wire w188018;

	wire w192018;

	wire w195018;

	wire w197018;

	wire w200018;

	wire w14019;

	wire w17019;

	wire w19019;

	wire w22019;

	wire w26019;

	wire w187019;

	wire w189019;

	wire w191019;

	wire w193019;

	wire w196019;

	wire w199019;

	wire w201019;

	wire w13020;

	wire w15020;

	wire w18020;

	wire w21020;

	wire w23020;

	wire w25020;

	wire w27020;

	wire w192020;

	wire w22021;

	wire w40021;
	torch #(1'b1) c40021 (.i_clk(tick), .i_in(), .o_out(w40021));
	wire w44021;
	torch #(1'b1) c44021 (.i_clk(tick), .i_in(), .o_out(w44021));
	wire w48021;
	torch #(1'b1) c48021 (.i_clk(tick), .i_in(), .o_out(w48021));
	wire w52021;
	torch #(1'b1) c52021 (.i_clk(tick), .i_in(), .o_out(w52021));
	wire w56021;
	torch #(1'b1) c56021 (.i_clk(tick), .i_in(), .o_out(w56021));
	wire w60021;
	torch #(1'b1) c60021 (.i_clk(tick), .i_in(), .o_out(w60021));
	wire w64021;
	torch #(1'b1) c64021 (.i_clk(tick), .i_in(), .o_out(w64021));
	wire w188021;

	wire w192021;

	wire w193021;

	wire w197021;

	wire w199021;

	wire w201021;

	wire w13022;

	wire w15022;

	wire w17022;

	wire w21022;

	wire w22022;

	wire w26022;

	wire w193023;

	wire w21024;

	wire w118026;

	wire w152026;

	wire w116027;
	repeater #(1, 1'b1, 0, 0) c116027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116027));
	wire w150027;
	repeater #(1, 1'b1, 0, 0) c150027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150027));
	wire w107028;
	repeater #(1, 1'b1, 0, 0) c107028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107028));
	wire w123028;
	repeater #(1, 1'b1, 0, 0) c123028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123028));
	wire w141028;
	repeater #(1, 1'b1, 0, 0) c141028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141028));
	wire w157028;
	repeater #(1, 1'b1, 0, 0) c157028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157028));
	wire w44029;
	repeater #(1, 1'b0, 0, 0) c44029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44029));
	wire w64029;
	repeater #(1, 1'b0, 0, 0) c64029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64029));
	wire w118029;

	wire w134029;

	wire w152029;

	wire w168029;

	wire w110030;

	wire w126030;

	wire w144030;

	wire w160030;

	wire w107031;

	wire w108031;

	wire w113031;

	wire w121031;

	wire w123031;

	wire w124031;

	wire w129031;

	wire w137031;

	wire w141031;

	wire w142031;

	wire w147031;

	wire w155031;

	wire w157031;

	wire w158031;

	wire w163031;

	wire w171031;

	wire w115033;

	wire w116033;

	wire w131033;

	wire w132033;

	wire w149033;

	wire w150033;

	wire w165033;

	wire w166033;

	wire w107035;

	wire w108035;

	wire w121035;

	wire w123035;

	wire w124035;

	wire w137035;

	wire w141035;

	wire w142035;

	wire w155035;

	wire w157035;

	wire w158035;

	wire w171035;

	wire w1036;

	wire w200036;
	repeater #(1, 1'b1, 0, 0) c200036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200036));
	wire w14037;
	repeater #(1, 1'b1, 0, 0) c14037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14037));
	wire w40037;
	torch #(1'b1) c40037 (.i_clk(tick), .i_in(), .o_out(w40037));
	wire w44037;
	torch #(1'b1) c44037 (.i_clk(tick), .i_in(), .o_out(w44037));
	wire w48037;
	torch #(1'b1) c48037 (.i_clk(tick), .i_in(), .o_out(w48037));
	wire w52037;
	torch #(1'b1) c52037 (.i_clk(tick), .i_in(), .o_out(w52037));
	wire w56037;
	torch #(1'b1) c56037 (.i_clk(tick), .i_in(), .o_out(w56037));
	wire w60037;
	torch #(1'b1) c60037 (.i_clk(tick), .i_in(), .o_out(w60037));
	wire w64037;
	torch #(1'b1) c64037 (.i_clk(tick), .i_in(), .o_out(w64037));
	wire w118037;
	torch #(1'b1) c118037 (.i_clk(tick), .i_in(), .o_out(w118037));
	wire w119037;

	wire w134037;
	torch #(1'b1) c134037 (.i_clk(tick), .i_in(), .o_out(w134037));
	wire w135037;

	wire w152037;
	torch #(1'b1) c152037 (.i_clk(tick), .i_in(), .o_out(w152037));
	wire w153037;

	wire w168037;
	torch #(1'b1) c168037 (.i_clk(tick), .i_in(), .o_out(w168037));
	wire w169037;

	wire w3038;

	wire w119038;

	wire w121038;

	wire w135038;

	wire w137038;

	wire w153038;

	wire w155038;

	wire w169038;

	wire w171038;

	wire w4039;

	wire w203039;
	repeater #(1, 1'b1, 0, 0) c203039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203039));
	wire w204039;

	wire w4040;
	repeater #(1, 1'b0, 0, 0) c4040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4040));
	wire w10040;

	wire w11040;
	repeater #(1, 1'b1, 0, 0) c11040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11040));
	wire w121040;

	wire w122040;

	wire w123040;

	wire w137040;

	wire w138040;

	wire w139040;

	wire w155040;

	wire w156040;

	wire w157040;

	wire w171040;

	wire w172040;

	wire w173040;

	wire w200040;

	wire w201040;

	wire w13041;

	wire w14041;

	wire w116041;

	wire w117041;

	wire w123041;

	wire w132041;

	wire w133041;

	wire w139041;

	wire w150041;

	wire w151041;

	wire w157041;

	wire w166041;

	wire w167041;

	wire w173041;

	wire w3042;

	wire w4042;

	wire w200042;
	repeater #(1, 1'b1, 0, 0) c200042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200042));
	wire w0043;

	wire w1043;
	repeater #(1, 1'b1, 0, 0) c1043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1043));
	wire w14043;
	repeater #(1, 1'b0, 0, 0) c14043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14043));
	wire w113043;
	torch #(1'b0) c113043 (.i_clk(tick), .i_in(), .o_out(w113043));
	wire w121043;
	repeater #(1, 1'b0, 0, 0) c121043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121043));
	wire w123043;
	torch #(1'b0) c123043 (.i_clk(tick), .i_in(), .o_out(w123043));
	wire w129043;
	torch #(1'b0) c129043 (.i_clk(tick), .i_in(), .o_out(w129043));
	wire w137043;
	repeater #(1, 1'b0, 0, 0) c137043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137043));
	wire w139043;
	torch #(1'b0) c139043 (.i_clk(tick), .i_in(), .o_out(w139043));
	wire w147043;
	torch #(1'b0) c147043 (.i_clk(tick), .i_in(), .o_out(w147043));
	wire w155043;
	repeater #(1, 1'b0, 0, 0) c155043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155043));
	wire w157043;
	torch #(1'b0) c157043 (.i_clk(tick), .i_in(), .o_out(w157043));
	wire w163043;
	torch #(1'b0) c163043 (.i_clk(tick), .i_in(), .o_out(w163043));
	wire w171043;
	repeater #(1, 1'b0, 0, 0) c171043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171043));
	wire w173043;
	torch #(1'b0) c173043 (.i_clk(tick), .i_in(), .o_out(w173043));
	wire w200043;

	wire w9044;

	wire w14044;

	wire w201044;

	wire w205044;
	repeater #(1, 1'b1, 0, 0) c205044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205044));
	wire w10045;
	repeater #(2, 1'b0, 0, 0) c10045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10045));
	wire w13045;

	wire w44045;
	repeater #(1, 1'b0, 0, 0) c44045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44045));
	wire w64045;
	repeater #(1, 1'b0, 0, 0) c64045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64045));
	wire w125045;
	repeater #(1, 1'b0, 0, 0) c125045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125045));
	wire w159045;
	repeater #(1, 1'b0, 0, 0) c159045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159045));
	wire w204045;
	assign outputs[53] = ();
	wire w122047;
	torch #(1'b1) c122047 (.i_clk(tick), .i_in(), .o_out(w122047));
	wire w138047;
	torch #(1'b1) c138047 (.i_clk(tick), .i_in(), .o_out(w138047));
	wire w156047;
	torch #(1'b1) c156047 (.i_clk(tick), .i_in(), .o_out(w156047));
	wire w172047;
	torch #(1'b1) c172047 (.i_clk(tick), .i_in(), .o_out(w172047));
	wire w114049;
	torch #(1'b1) c114049 (.i_clk(tick), .i_in(), .o_out(w114049));
	wire w130049;
	torch #(1'b1) c130049 (.i_clk(tick), .i_in(), .o_out(w130049));
	wire w148049;
	torch #(1'b1) c148049 (.i_clk(tick), .i_in(), .o_out(w148049));
	wire w164049;
	torch #(1'b1) c164049 (.i_clk(tick), .i_in(), .o_out(w164049));
	wire w121050;
	repeater #(2, 1'b0, 0, 0) c121050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121050));
	wire w137050;
	repeater #(1, 1'b0, 0, 0) c137050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137050));
	wire w155050;
	repeater #(2, 1'b0, 0, 0) c155050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155050));
	wire w171050;
	repeater #(1, 1'b0, 0, 0) c171050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171050));
	wire w115051;
	repeater #(2, 1'b0, 0, 0) c115051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115051));
	wire w131051;
	repeater #(1, 1'b0, 0, 0) c131051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131051));
	wire w149051;
	repeater #(2, 1'b0, 0, 0) c149051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149051));
	wire w165051;
	repeater #(1, 1'b0, 0, 0) c165051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165051));
	wire w40053;
	torch #(1'b1) c40053 (.i_clk(tick), .i_in(), .o_out(w40053));
	wire w44053;
	torch #(1'b1) c44053 (.i_clk(tick), .i_in(), .o_out(w44053));
	wire w48053;
	torch #(1'b1) c48053 (.i_clk(tick), .i_in(), .o_out(w48053));
	wire w52053;
	torch #(1'b1) c52053 (.i_clk(tick), .i_in(), .o_out(w52053));
	wire w56053;
	torch #(1'b1) c56053 (.i_clk(tick), .i_in(), .o_out(w56053));
	wire w60053;
	torch #(1'b1) c60053 (.i_clk(tick), .i_in(), .o_out(w60053));
	wire w64053;
	torch #(1'b1) c64053 (.i_clk(tick), .i_in(), .o_out(w64053));
	wire w125053;
	repeater #(1, 1'b0, 0, 0) c125053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125053));
	wire w159053;
	repeater #(1, 1'b0, 0, 0) c159053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159053));
	wire w127054;
	repeater #(1, 1'b0, 0, 0) c127054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127054));
	wire w161054;
	repeater #(1, 1'b0, 0, 0) c161054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161054));
	wire w44061;
	repeater #(1, 1'b0, 0, 0) c44061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44061));
	wire w64061;
	repeater #(1, 1'b0, 0, 0) c64061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64061));
	wire w2068;

	wire w3068;
	repeater #(1, 1'b0, 0, 0) c3068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3068));
	wire w4069;
	repeater #(1, 1'b0, 0, 0) c4069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4069));
	wire w7069;
	repeater #(2, 1'b0, 0, 0) c7069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7069));
	wire w40069;
	torch #(1'b1) c40069 (.i_clk(tick), .i_in(), .o_out(w40069));
	wire w44069;
	torch #(1'b1) c44069 (.i_clk(tick), .i_in(), .o_out(w44069));
	wire w48069;
	torch #(1'b1) c48069 (.i_clk(tick), .i_in(), .o_out(w48069));
	wire w52069;
	torch #(1'b1) c52069 (.i_clk(tick), .i_in(), .o_out(w52069));
	wire w56069;
	torch #(1'b1) c56069 (.i_clk(tick), .i_in(), .o_out(w56069));
	wire w60069;
	torch #(1'b1) c60069 (.i_clk(tick), .i_in(), .o_out(w60069));
	wire w64069;
	torch #(1'b1) c64069 (.i_clk(tick), .i_in(), .o_out(w64069));
	wire w207069;
	repeater #(1, 1'b0, 0, 0) c207069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207069));
	wire w12070;
	repeater #(2, 1'b0, 0, 0) c12070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12070));
	wire w206070;
	assign outputs[54] = ();
	wire w1071;

	wire w10071;

	wire w1072;

	wire w10072;

	wire w207072;
	repeater #(1, 1'b0, 0, 0) c207072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207072));
	wire w12073;
	repeater #(1, 1'b0, 0, 0) c12073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12073));
	wire w44077;
	repeater #(1, 1'b0, 0, 0) c44077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44077));
	wire w64077;
	repeater #(1, 1'b0, 0, 0) c64077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64077));
	wire w40085;
	torch #(1'b1) c40085 (.i_clk(tick), .i_in(), .o_out(w40085));
	wire w44085;
	torch #(1'b1) c44085 (.i_clk(tick), .i_in(), .o_out(w44085));
	wire w48085;
	torch #(1'b1) c48085 (.i_clk(tick), .i_in(), .o_out(w48085));
	wire w52085;
	torch #(1'b1) c52085 (.i_clk(tick), .i_in(), .o_out(w52085));
	wire w56085;
	torch #(1'b1) c56085 (.i_clk(tick), .i_in(), .o_out(w56085));
	wire w60085;
	torch #(1'b1) c60085 (.i_clk(tick), .i_in(), .o_out(w60085));
	wire w64085;
	torch #(1'b1) c64085 (.i_clk(tick), .i_in(), .o_out(w64085));
	wire w41098;
	torch #(1'b1) c41098 (.i_clk(tick), .i_in(), .o_out(w41098));
	wire w45098;
	torch #(1'b1) c45098 (.i_clk(tick), .i_in(), .o_out(w45098));
	wire w49098;
	torch #(1'b1) c49098 (.i_clk(tick), .i_in(), .o_out(w49098));
	wire w53098;
	torch #(1'b1) c53098 (.i_clk(tick), .i_in(), .o_out(w53098));
	wire w57098;
	torch #(1'b1) c57098 (.i_clk(tick), .i_in(), .o_out(w57098));
	wire w61098;
	torch #(1'b1) c61098 (.i_clk(tick), .i_in(), .o_out(w61098));
	wire w65098;
	torch #(1'b1) c65098 (.i_clk(tick), .i_in(), .o_out(w65098));
	wire w410102;
	torch #(1'b1) c410102 (.i_clk(tick), .i_in(), .o_out(w410102));
	wire w450102;
	torch #(1'b1) c450102 (.i_clk(tick), .i_in(), .o_out(w450102));
	wire w490102;
	torch #(1'b1) c490102 (.i_clk(tick), .i_in(), .o_out(w490102));
	wire w530102;
	torch #(1'b0) c530102 (.i_clk(tick), .i_in(), .o_out(w530102));
	wire w570102;
	torch #(1'b1) c570102 (.i_clk(tick), .i_in(), .o_out(w570102));
	wire w610102;
	torch #(1'b1) c610102 (.i_clk(tick), .i_in(), .o_out(w610102));
	wire w650102;
	torch #(1'b1) c650102 (.i_clk(tick), .i_in(), .o_out(w650102));
	wire w400110;
	torch #(1'b1) c400110 (.i_clk(tick), .i_in(), .o_out(w400110));
	wire w440110;
	torch #(1'b1) c440110 (.i_clk(tick), .i_in(), .o_out(w440110));
	wire w480110;
	torch #(1'b1) c480110 (.i_clk(tick), .i_in(), .o_out(w480110));
	wire w520110;
	torch #(1'b1) c520110 (.i_clk(tick), .i_in(), .o_out(w520110));
	wire w560110;
	torch #(1'b1) c560110 (.i_clk(tick), .i_in(), .o_out(w560110));
	wire w600110;
	torch #(1'b1) c600110 (.i_clk(tick), .i_in(), .o_out(w600110));
	wire w640110;
	torch #(1'b1) c640110 (.i_clk(tick), .i_in(), .o_out(w640110));
	wire w390120;
	repeater #(1, 1'b0, 0, 0) c390120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390120));
	wire w430120;
	repeater #(1, 1'b0, 0, 0) c430120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w430120));
	wire w470120;
	repeater #(1, 1'b0, 0, 0) c470120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470120));
	wire w510120;
	repeater #(1, 1'b0, 0, 0) c510120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w510120));
	wire w550120;
	repeater #(1, 1'b0, 0, 0) c550120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550120));
	wire w590120;
	repeater #(1, 1'b0, 0, 0) c590120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w590120));
	wire w630120;
	repeater #(1, 1'b0, 0, 0) c630120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630120));
	wire w410143;
	repeater #(1, 1'b0, 0, 0) c410143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w410143));
	wire w450143;
	repeater #(1, 1'b0, 0, 0) c450143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w450143));
	wire w490143;
	repeater #(1, 1'b0, 0, 0) c490143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w490143));
	wire w530143;
	repeater #(1, 1'b0, 0, 0) c530143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530143));
	wire w570143;
	repeater #(1, 1'b0, 0, 0) c570143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570143));
	wire w610143;
	repeater #(1, 1'b0, 0, 0) c610143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w610143));
	wire w650143;
	repeater #(1, 1'b0, 0, 0) c650143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650143));
	wire w410146;
	torch #(1'b1) c410146 (.i_clk(tick), .i_in(), .o_out(w410146));
	wire w450146;
	torch #(1'b1) c450146 (.i_clk(tick), .i_in(), .o_out(w450146));
	wire w490146;
	torch #(1'b1) c490146 (.i_clk(tick), .i_in(), .o_out(w490146));
	wire w530146;
	torch #(1'b1) c530146 (.i_clk(tick), .i_in(), .o_out(w530146));
	wire w570146;
	torch #(1'b1) c570146 (.i_clk(tick), .i_in(), .o_out(w570146));
	wire w610146;
	torch #(1'b1) c610146 (.i_clk(tick), .i_in(), .o_out(w610146));
	wire w650146;
	torch #(1'b1) c650146 (.i_clk(tick), .i_in(), .o_out(w650146));
	wire w520149;
	repeater #(1, 1'b0, 0, 0) c520149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520149));
	wire w540149;
	repeater #(1, 1'b1, 0, 0) c540149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540149));
	wire w560149;
	repeater #(1, 1'b1, 0, 0) c560149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560149));
	wire w580149;
	repeater #(1, 1'b1, 0, 0) c580149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580149));
	wire w600149;
	repeater #(1, 1'b1, 0, 0) c600149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600149));
	wire w620149;
	repeater #(1, 1'b1, 0, 0) c620149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620149));
	wire w640149;
	repeater #(1, 1'b1, 0, 0) c640149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640149));
	wire w660149;
	repeater #(1, 1'b1, 0, 0) c660149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660149));
	wire w500151;
	repeater #(1, 1'b1, 0, 0) c500151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500151));
	wire w480153;
	repeater #(1, 1'b1, 0, 0) c480153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480153));
	wire w460155;
	repeater #(1, 1'b1, 0, 0) c460155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460155));
	wire w440157;
	repeater #(1, 1'b1, 0, 0) c440157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440157));
	wire w420159;
	repeater #(1, 1'b1, 0, 0) c420159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420159));
	wire w400161;
	repeater #(1, 1'b1, 0, 0) c400161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400161));
	wire w1380166;
	torch #(1'b1) c1380166 (.i_clk(tick), .i_in(), .o_out(w1380166));
	wire w1720166;
	repeater #(1, 1'b1, 0, 0) c1720166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1720166));
	wire w2060166;
	torch #(1'b1) c2060166 (.i_clk(tick), .i_in(), .o_out(w2060166));
	wire w320167;
	repeater #(1, 1'b1, 0, 0) c320167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320167));
	wire w1360168;
	repeater #(1, 1'b1, 0, 0) c1360168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1360168));
	wire w1700168;
	repeater #(1, 1'b1, 0, 0) c1700168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1700168));
	wire w2040168;
	repeater #(1, 1'b1, 0, 0) c2040168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040168));
	wire w300169;
	repeater #(1, 1'b1, 0, 0) c300169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300169));
	wire w660170;
	repeater #(1, 1'b1, 0, 0) c660170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660170));
	wire w1340170;
	torch #(1'b1) c1340170 (.i_clk(tick), .i_in(), .o_out(w1340170));
	wire w1680170;
	repeater #(1, 1'b1, 0, 0) c1680170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1680170));
	wire w2020170;
	torch #(1'b1) c2020170 (.i_clk(tick), .i_in(), .o_out(w2020170));
	wire w280171;
	repeater #(1, 1'b1, 0, 0) c280171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280171));
	wire w640172;
	repeater #(1, 1'b1, 0, 0) c640172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640172));
	wire w1320172;
	repeater #(1, 1'b1, 0, 0) c1320172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1320172));
	wire w1660172;
	repeater #(1, 1'b1, 0, 0) c1660172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1660172));
	wire w2000172;
	repeater #(1, 1'b1, 0, 0) c2000172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2000172));
	wire w260173;
	repeater #(1, 1'b1, 0, 0) c260173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260173));
	wire w620174;
	repeater #(1, 1'b1, 0, 0) c620174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620174));
	wire w1300174;
	torch #(1'b1) c1300174 (.i_clk(tick), .i_in(), .o_out(w1300174));
	wire w1640174;
	repeater #(1, 1'b1, 0, 0) c1640174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640174));
	wire w1980174;
	torch #(1'b1) c1980174 (.i_clk(tick), .i_in(), .o_out(w1980174));
	wire w240175;
	repeater #(1, 1'b1, 0, 0) c240175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240175));
	wire w600176;
	repeater #(1, 1'b1, 0, 0) c600176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600176));
	wire w1280176;
	repeater #(1, 1'b1, 0, 0) c1280176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1280176));
	wire w1620176;
	repeater #(1, 1'b1, 0, 0) c1620176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620176));
	wire w1960176;
	repeater #(1, 1'b1, 0, 0) c1960176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1960176));
	wire w220177;
	repeater #(1, 1'b1, 0, 0) c220177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220177));
	wire w1120177;
	repeater #(1, 1'b1, 0, 0) c1120177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1120177));
	wire w1140177;
	torch #(1'b1) c1140177 (.i_clk(tick), .i_in(), .o_out(w1140177));
	wire w1160177;
	repeater #(1, 1'b1, 0, 0) c1160177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1160177));
	wire w1180177;
	torch #(1'b1) c1180177 (.i_clk(tick), .i_in(), .o_out(w1180177));
	wire w1200177;
	repeater #(1, 1'b1, 0, 0) c1200177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1200177));
	wire w1220177;
	torch #(1'b1) c1220177 (.i_clk(tick), .i_in(), .o_out(w1220177));
	wire w1240177;
	repeater #(1, 1'b0, 0, 0) c1240177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240177));
	wire w1260177;
	torch #(1'b1) c1260177 (.i_clk(tick), .i_in(), .o_out(w1260177));
	wire w1460177;
	repeater #(1, 1'b1, 0, 0) c1460177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460177));
	wire w1480177;
	repeater #(1, 1'b1, 0, 0) c1480177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1480177));
	wire w1500177;
	repeater #(1, 1'b1, 0, 0) c1500177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500177));
	wire w1520177;
	repeater #(1, 1'b1, 0, 0) c1520177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520177));
	wire w1540177;
	repeater #(1, 1'b1, 0, 0) c1540177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540177));
	wire w1560177;
	repeater #(1, 1'b1, 0, 0) c1560177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560177));
	wire w1580177;
	repeater #(1, 1'b0, 0, 0) c1580177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580177));
	wire w1600177;
	repeater #(1, 1'b1, 0, 0) c1600177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1600177));
	wire w1820177;
	torch #(1'b1) c1820177 (.i_clk(tick), .i_in(), .o_out(w1820177));
	wire w1860177;
	torch #(1'b1) c1860177 (.i_clk(tick), .i_in(), .o_out(w1860177));
	wire w1900177;
	torch #(1'b1) c1900177 (.i_clk(tick), .i_in(), .o_out(w1900177));
	wire w1940177;
	torch #(1'b1) c1940177 (.i_clk(tick), .i_in(), .o_out(w1940177));
	wire w60178;
	repeater #(1, 1'b1, 0, 0) c60178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60178));
	wire w80178;
	repeater #(1, 1'b1, 0, 0) c80178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80178));
	wire w100178;
	repeater #(1, 1'b1, 0, 0) c100178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100178));
	wire w120178;
	repeater #(1, 1'b1, 0, 0) c120178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120178));
	wire w140178;
	repeater #(1, 1'b1, 0, 0) c140178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140178));
	wire w160178;
	repeater #(1, 1'b1, 0, 0) c160178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160178));
	wire w180178;
	repeater #(1, 1'b0, 0, 0) c180178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180178));
	wire w200178;
	repeater #(1, 1'b1, 0, 0) c200178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200178));
	wire w580178;
	repeater #(1, 1'b1, 0, 0) c580178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580178));
	wire w1810178;
	repeater #(1, 1'b1, 0, 0) c1810178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810178));
	wire w1850178;
	repeater #(1, 1'b1, 0, 0) c1850178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850178));
	wire w1890178;
	repeater #(1, 1'b1, 0, 0) c1890178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1890178));
	wire w1930178;
	repeater #(1, 1'b0, 0, 0) c1930178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1930178));
	wire w4410;
	repeater #(1, 1'b1, 0, 0) c4410 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4410));
	wire w4610;
	repeater #(1, 1'b1, 0, 0) c4610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4610));
	wire w4810;
	repeater #(1, 1'b1, 0, 0) c4810 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4810));
	wire w5010;
	repeater #(1, 1'b1, 0, 0) c5010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5010));
	wire w5210;
	repeater #(1, 1'b0, 0, 0) c5210 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5210));
	wire w5410;
	repeater #(1, 1'b1, 0, 0) c5410 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5410));
	wire w5610;
	repeater #(1, 1'b1, 0, 0) c5610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5610));
	wire w18211;
	torch #(1'b1) c18211 (.i_clk(tick), .i_in(), .o_out(w18211));
	wire w18611;
	torch #(1'b1) c18611 (.i_clk(tick), .i_in(), .o_out(w18611));
	wire w19011;
	torch #(1'b1) c19011 (.i_clk(tick), .i_in(), .o_out(w19011));
	wire w19411;
	torch #(1'b0) c19411 (.i_clk(tick), .i_in(), .o_out(w19411));
	wire w19811;
	torch #(1'b1) c19811 (.i_clk(tick), .i_in(), .o_out(w19811));
	wire w20211;
	torch #(1'b1) c20211 (.i_clk(tick), .i_in(), .o_out(w20211));
	wire w20611;
	torch #(1'b1) c20611 (.i_clk(tick), .i_in(), .o_out(w20611));
	wire w812;
	torch #(1'b1) c812 (.i_clk(tick), .i_in(), .o_out(w812));
	wire w1212;
	torch #(1'b1) c1212 (.i_clk(tick), .i_in(), .o_out(w1212));
	wire w1612;
	torch #(1'b1) c1612 (.i_clk(tick), .i_in(), .o_out(w1612));
	wire w2012;
	torch #(1'b1) c2012 (.i_clk(tick), .i_in(), .o_out(w2012));
	wire w2412;
	torch #(1'b1) c2412 (.i_clk(tick), .i_in(), .o_out(w2412));
	wire w2812;
	torch #(1'b1) c2812 (.i_clk(tick), .i_in(), .o_out(w2812));
	wire w3212;
	torch #(1'b1) c3212 (.i_clk(tick), .i_in(), .o_out(w3212));
	wire w11212;
	repeater #(2, 1'b1, 0, 0) c11212 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11212));
	wire w11612;
	repeater #(2, 1'b1, 0, 0) c11612 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11612));
	wire w12012;
	repeater #(2, 1'b1, 0, 0) c12012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12012));
	wire w13612;
	repeater #(2, 1'b0, 0, 0) c13612 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13612));
	wire w14612;
	repeater #(2, 1'b1, 0, 0) c14612 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14612));
	wire w15012;
	repeater #(2, 1'b1, 0, 0) c15012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15012));
	wire w15412;
	repeater #(2, 1'b1, 0, 0) c15412 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15412));
	wire w17012;
	repeater #(2, 1'b0, 0, 0) c17012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17012));
	wire w18713;
	torch #(1'b1) c18713 (.i_clk(tick), .i_in(), .o_out(w18713));
	wire w19113;
	torch #(1'b1) c19113 (.i_clk(tick), .i_in(), .o_out(w19113));
	wire w19513;
	torch #(1'b1) c19513 (.i_clk(tick), .i_in(), .o_out(w19513));
	wire w19913;
	torch #(1'b1) c19913 (.i_clk(tick), .i_in(), .o_out(w19913));
	wire w1514;
	torch #(1'b0) c1514 (.i_clk(tick), .i_in(), .o_out(w1514));
	wire w1914;
	torch #(1'b0) c1914 (.i_clk(tick), .i_in(), .o_out(w1914));
	wire w2314;
	torch #(1'b0) c2314 (.i_clk(tick), .i_in(), .o_out(w2314));
	wire w2714;
	torch #(1'b0) c2714 (.i_clk(tick), .i_in(), .o_out(w2714));
	wire w11214;
	torch #(1'b1) c11214 (.i_clk(tick), .i_in(), .o_out(w11214));
	wire w12214;
	repeater #(1, 1'b1, 0, 0) c12214 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12214));
	wire w12814;
	torch #(1'b1) c12814 (.i_clk(tick), .i_in(), .o_out(w12814));
	wire w13814;
	repeater #(1, 1'b0, 0, 0) c13814 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13814));
	wire w14614;
	torch #(1'b1) c14614 (.i_clk(tick), .i_in(), .o_out(w14614));
	wire w15614;
	repeater #(1, 1'b1, 0, 0) c15614 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15614));
	wire w16214;
	torch #(1'b1) c16214 (.i_clk(tick), .i_in(), .o_out(w16214));
	wire w17214;
	repeater #(1, 1'b1, 0, 0) c17214 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17214));
	wire w12917;
	repeater #(1, 1'b1, 0, 0) c12917 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12917));
	wire w16317;
	repeater #(1, 1'b1, 0, 0) c16317 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16317));
	wire w12218;
	repeater #(1, 1'b1, 0, 0) c12218 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12218));
	wire w13818;
	repeater #(1, 1'b0, 0, 0) c13818 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13818));
	wire w15618;
	repeater #(1, 1'b1, 0, 0) c15618 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15618));
	wire w17218;
	repeater #(1, 1'b1, 0, 0) c17218 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17218));
	wire w11119;

	wire w12719;

	wire w14519;

	wire w16119;

	wire w42110;
	repeater #(1, 1'b1, 0, 0) c42110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42110));
	wire w46110;
	repeater #(1, 1'b1, 0, 0) c46110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46110));
	wire w50110;
	repeater #(1, 1'b1, 0, 0) c50110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50110));
	wire w54110;
	repeater #(1, 1'b0, 0, 0) c54110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54110));
	wire w58110;
	repeater #(1, 1'b1, 0, 0) c58110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58110));
	wire w62110;
	repeater #(1, 1'b1, 0, 0) c62110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62110));
	wire w66110;
	repeater #(1, 1'b1, 0, 0) c66110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66110));
	wire w119110;

	wire w135110;

	wire w153110;

	wire w169110;

	wire w116111;

	wire w121111;

	wire w122111;

	wire w132111;

	wire w137111;

	wire w138111;

	wire w150111;

	wire w155111;

	wire w156111;

	wire w166111;

	wire w171111;

	wire w172111;

	wire w114113;

	wire w130113;

	wire w148113;

	wire w164113;

	wire w44114;

	wire w69114;
	repeater #(1, 1'b0, 0, 0) c69114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69114));
	wire w120114;

	wire w121114;

	wire w136114;

	wire w137114;

	wire w154114;

	wire w155114;

	wire w170114;

	wire w171114;

	wire w64115;

	wire w130115;

	wire w134115;

	wire w164115;

	wire w168115;

	wire w39116;
	repeater #(1, 1'b0, 0, 0) c39116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39116));
	wire w48119;
	torch #(1'b1) c48119 (.i_clk(tick), .i_in(), .o_out(w48119));
	wire w52119;
	torch #(1'b1) c52119 (.i_clk(tick), .i_in(), .o_out(w52119));
	wire w56119;
	torch #(1'b1) c56119 (.i_clk(tick), .i_in(), .o_out(w56119));
	wire w60119;
	torch #(1'b1) c60119 (.i_clk(tick), .i_in(), .o_out(w60119));
	wire w111119;

	wire w112119;

	wire w115119;

	wire w116119;

	wire w119119;

	wire w120119;

	wire w123119;

	wire w124119;

	wire w127119;

	wire w128119;

	wire w131119;

	wire w132119;

	wire w135119;

	wire w136119;

	wire w145119;

	wire w146119;

	wire w149119;

	wire w150119;

	wire w153119;

	wire w154119;

	wire w157119;

	wire w158119;

	wire w161119;

	wire w162119;

	wire w165119;

	wire w166119;

	wire w169119;

	wire w170119;

	wire w112121;

	wire w116121;

	wire w120121;

	wire w124121;

	wire w128121;

	wire w132121;

	wire w136121;

	wire w146121;

	wire w150121;

	wire w154121;

	wire w158121;

	wire w162121;

	wire w166121;

	wire w170121;

	wire w41123;
	torch #(1'b0) c41123 (.i_clk(tick), .i_in(), .o_out(w41123));
	wire w45123;
	torch #(1'b0) c45123 (.i_clk(tick), .i_in(), .o_out(w45123));
	wire w49123;
	torch #(1'b0) c49123 (.i_clk(tick), .i_in(), .o_out(w49123));
	wire w53123;
	torch #(1'b1) c53123 (.i_clk(tick), .i_in(), .o_out(w53123));
	wire w57123;
	torch #(1'b0) c57123 (.i_clk(tick), .i_in(), .o_out(w57123));
	wire w61123;
	torch #(1'b0) c61123 (.i_clk(tick), .i_in(), .o_out(w61123));
	wire w65123;
	torch #(1'b0) c65123 (.i_clk(tick), .i_in(), .o_out(w65123));
	wire w110124;

	wire w114124;

	wire w118124;

	wire w122124;

	wire w144124;

	wire w148124;

	wire w152124;

	wire w156124;

	wire w190124;

	wire w191124;
	repeater #(2, 1'b1, 0, 0) c191124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191124));
	wire w23125;
	repeater #(2, 1'b1, 0, 0) c23125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23125));
	wire w24125;

	wire w42125;
	torch #(1'b1) c42125 (.i_clk(tick), .i_in(), .o_out(w42125));
	wire w46125;
	torch #(1'b1) c46125 (.i_clk(tick), .i_in(), .o_out(w46125));
	wire w50125;
	torch #(1'b1) c50125 (.i_clk(tick), .i_in(), .o_out(w50125));
	wire w54125;
	torch #(1'b1) c54125 (.i_clk(tick), .i_in(), .o_out(w54125));
	wire w58125;
	torch #(1'b1) c58125 (.i_clk(tick), .i_in(), .o_out(w58125));
	wire w62125;
	torch #(1'b1) c62125 (.i_clk(tick), .i_in(), .o_out(w62125));
	wire w66125;
	torch #(1'b1) c66125 (.i_clk(tick), .i_in(), .o_out(w66125));
	wire w183125;
	repeater #(1, 1'b1, 0, 0) c183125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183125));
	wire w188125;
	repeater #(1, 1'b1, 0, 0) c188125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188125));
	wire w193125;
	repeater #(1, 1'b1, 0, 0) c193125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193125));
	wire w21126;
	repeater #(1, 1'b1, 0, 0) c21126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21126));
	wire w26126;
	repeater #(1, 1'b1, 0, 0) c26126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26126));
	wire w31126;
	repeater #(1, 1'b1, 0, 0) c31126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31126));
	wire w122126;

	wire w156126;

	wire w182126;

	wire w183126;
	repeater #(1, 1'b1, 0, 0) c183126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183126));
	wire w187126;

	wire w188126;
	repeater #(1, 1'b1, 0, 0) c188126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188126));
	wire w192126;

	wire w193126;
	repeater #(1, 1'b1, 0, 0) c193126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193126));
	wire w21127;
	repeater #(1, 1'b1, 0, 0) c21127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21127));
	wire w22127;

	wire w26127;
	repeater #(1, 1'b1, 0, 0) c26127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26127));
	wire w27127;

	wire w31127;
	repeater #(1, 1'b1, 0, 0) c31127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31127));
	wire w32127;

	wire w120127;
	repeater #(1, 1'b1, 0, 0) c120127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120127));
	wire w154127;
	repeater #(1, 1'b1, 0, 0) c154127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154127));
	wire w111128;
	repeater #(1, 1'b1, 0, 0) c111128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111128));
	wire w127128;
	repeater #(1, 1'b1, 0, 0) c127128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127128));
	wire w145128;
	repeater #(1, 1'b1, 0, 0) c145128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145128));
	wire w161128;
	repeater #(1, 1'b1, 0, 0) c161128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161128));
	wire w122129;

	wire w156129;

	wire w183129;
	repeater #(1, 1'b1, 0, 0) c183129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183129));
	wire w188129;
	repeater #(1, 1'b1, 0, 0) c188129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188129));
	wire w193129;
	repeater #(1, 1'b1, 0, 0) c193129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193129));
	wire w21130;
	repeater #(1, 1'b1, 0, 0) c21130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21130));
	wire w26130;
	repeater #(1, 1'b1, 0, 0) c26130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26130));
	wire w31130;
	repeater #(1, 1'b1, 0, 0) c31130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31130));
	wire w44130;

	wire w69130;
	repeater #(1, 1'b0, 0, 0) c69130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69130));
	wire w114130;

	wire w148130;

	wire w182130;

	wire w183130;
	repeater #(1, 1'b0, 0, 0) c183130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183130));
	wire w187130;

	wire w188130;
	repeater #(1, 1'b0, 0, 0) c188130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188130));
	wire w192130;

	wire w193130;
	repeater #(1, 1'b1, 0, 0) c193130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193130));
	wire w21131;
	repeater #(1, 1'b1, 0, 0) c21131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21131));
	wire w22131;

	wire w26131;
	repeater #(1, 1'b0, 0, 0) c26131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26131));
	wire w27131;

	wire w31131;
	repeater #(1, 1'b1, 0, 0) c31131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31131));
	wire w32131;

	wire w64131;

	wire w111131;

	wire w112131;

	wire w117131;

	wire w125131;

	wire w127131;

	wire w128131;

	wire w145131;

	wire w146131;

	wire w151131;

	wire w159131;

	wire w161131;

	wire w162131;

	wire w39132;
	repeater #(1, 1'b0, 0, 0) c39132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39132));
	wire w119133;

	wire w120133;

	wire w153133;

	wire w154133;

	wire w183133;
	repeater #(1, 1'b0, 0, 0) c183133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183133));
	wire w188133;
	repeater #(1, 1'b0, 0, 0) c188133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188133));
	wire w193133;
	repeater #(1, 1'b0, 0, 0) c193133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193133));
	wire w202133;
	repeater #(1, 1'b0, 0, 0) c202133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202133));
	wire w12134;
	repeater #(1, 1'b0, 0, 0) c12134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12134));
	wire w21134;
	repeater #(1, 1'b1, 0, 0) c21134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21134));
	wire w26134;
	repeater #(1, 1'b0, 0, 0) c26134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26134));
	wire w31134;
	repeater #(1, 1'b0, 0, 0) c31134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31134));
	wire w182134;

	wire w183134;
	repeater #(1, 1'b0, 0, 0) c183134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183134));
	wire w187134;

	wire w188134;
	repeater #(1, 1'b0, 0, 0) c188134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188134));
	wire w192134;

	wire w193134;
	repeater #(1, 1'b0, 0, 0) c193134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193134));
	wire w21135;
	repeater #(1, 1'b1, 0, 0) c21135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21135));
	wire w22135;

	wire w26135;
	repeater #(1, 1'b0, 0, 0) c26135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26135));
	wire w27135;

	wire w31135;
	repeater #(1, 1'b0, 0, 0) c31135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31135));
	wire w32135;

	wire w48135;
	torch #(1'b1) c48135 (.i_clk(tick), .i_in(), .o_out(w48135));
	wire w52135;
	torch #(1'b1) c52135 (.i_clk(tick), .i_in(), .o_out(w52135));
	wire w56135;
	torch #(1'b1) c56135 (.i_clk(tick), .i_in(), .o_out(w56135));
	wire w60135;
	torch #(1'b1) c60135 (.i_clk(tick), .i_in(), .o_out(w60135));
	wire w111135;

	wire w112135;

	wire w125135;

	wire w127135;

	wire w128135;

	wire w145135;

	wire w146135;

	wire w159135;

	wire w161135;

	wire w162135;

	wire w1137;
	repeater #(1, 1'b1, 0, 0) c1137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1137));
	wire w122137;
	torch #(1'b1) c122137 (.i_clk(tick), .i_in(), .o_out(w122137));
	wire w123137;

	wire w156137;
	torch #(1'b1) c156137 (.i_clk(tick), .i_in(), .o_out(w156137));
	wire w157137;

	wire w123138;

	wire w125138;

	wire w157138;

	wire w159138;

	wire w181138;
	repeater #(1, 1'b1, 0, 0) c181138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181138));
	wire w5139;

	wire w33139;
	repeater #(1, 1'b0, 0, 0) c33139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33139));
	wire w41139;
	torch #(1'b0) c41139 (.i_clk(tick), .i_in(), .o_out(w41139));
	wire w45139;
	torch #(1'b0) c45139 (.i_clk(tick), .i_in(), .o_out(w45139));
	wire w49139;
	torch #(1'b0) c49139 (.i_clk(tick), .i_in(), .o_out(w49139));
	wire w53139;
	torch #(1'b0) c53139 (.i_clk(tick), .i_in(), .o_out(w53139));
	wire w57139;
	torch #(1'b0) c57139 (.i_clk(tick), .i_in(), .o_out(w57139));
	wire w61139;
	torch #(1'b0) c61139 (.i_clk(tick), .i_in(), .o_out(w61139));
	wire w65139;
	torch #(1'b0) c65139 (.i_clk(tick), .i_in(), .o_out(w65139));
	wire w2140;

	wire w125140;

	wire w126140;

	wire w127140;

	wire w159140;

	wire w160140;

	wire w161140;

	wire w195140;
	repeater #(1, 1'b0, 0, 0) c195140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195140));
	wire w1141;

	wire w3141;
	repeater #(2, 1'b0, 0, 0) c3141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3141));
	wire w6141;
	repeater #(2, 1'b1, 0, 0) c6141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6141));
	wire w19141;
	repeater #(1, 1'b1, 0, 0) c19141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19141));
	wire w42141;
	torch #(1'b1) c42141 (.i_clk(tick), .i_in(), .o_out(w42141));
	wire w46141;
	torch #(1'b1) c46141 (.i_clk(tick), .i_in(), .o_out(w46141));
	wire w50141;
	torch #(1'b1) c50141 (.i_clk(tick), .i_in(), .o_out(w50141));
	wire w54141;
	torch #(1'b1) c54141 (.i_clk(tick), .i_in(), .o_out(w54141));
	wire w58141;
	torch #(1'b1) c58141 (.i_clk(tick), .i_in(), .o_out(w58141));
	wire w62141;
	torch #(1'b1) c62141 (.i_clk(tick), .i_in(), .o_out(w62141));
	wire w66141;
	torch #(1'b1) c66141 (.i_clk(tick), .i_in(), .o_out(w66141));
	wire w120141;

	wire w121141;

	wire w127141;

	wire w136141;

	wire w137141;

	wire w154141;

	wire w155141;

	wire w161141;

	wire w170141;

	wire w171141;

	wire w192141;

	wire w198141;
	repeater #(2, 1'b1, 0, 0) c198141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198141));
	wire w201141;
	repeater #(2, 1'b0, 0, 0) c201141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201141));
	wire w203141;

	wire w11142;

	wire w13142;
	repeater #(2, 1'b0, 0, 0) c13142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13142));
	wire w16142;
	repeater #(2, 1'b1, 0, 0) c16142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16142));
	wire w22142;

	wire w191142;
	repeater #(2, 1'b0, 0, 0) c191142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191142));
	wire w202142;

	wire w12143;

	wire w23143;
	repeater #(2, 1'b1, 0, 0) c23143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23143));
	wire w117143;
	torch #(1'b0) c117143 (.i_clk(tick), .i_in(), .o_out(w117143));
	wire w125143;
	repeater #(1, 1'b0, 0, 0) c125143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125143));
	wire w127143;
	torch #(1'b0) c127143 (.i_clk(tick), .i_in(), .o_out(w127143));
	wire w133143;
	torch #(1'b0) c133143 (.i_clk(tick), .i_in(), .o_out(w133143));
	wire w151143;
	torch #(1'b0) c151143 (.i_clk(tick), .i_in(), .o_out(w151143));
	wire w159143;
	repeater #(1, 1'b0, 0, 0) c159143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159143));
	wire w161143;
	torch #(1'b0) c161143 (.i_clk(tick), .i_in(), .o_out(w161143));
	wire w167143;
	torch #(1'b0) c167143 (.i_clk(tick), .i_in(), .o_out(w167143));
	wire w199143;

	wire w15144;

	wire w113145;
	repeater #(1, 1'b1, 0, 0) c113145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113145));
	wire w129145;
	repeater #(1, 1'b1, 0, 0) c129145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w129145));
	wire w147145;
	repeater #(1, 1'b1, 0, 0) c147145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147145));
	wire w163145;
	repeater #(1, 1'b1, 0, 0) c163145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163145));
	wire w9146;
	assign outputs[55] = ();
	wire w44146;

	wire w69146;
	repeater #(1, 1'b0, 0, 0) c69146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69146));
	wire w64147;

	wire w126147;
	torch #(1'b1) c126147 (.i_clk(tick), .i_in(), .o_out(w126147));
	wire w160147;
	torch #(1'b1) c160147 (.i_clk(tick), .i_in(), .o_out(w160147));
	wire w39148;
	repeater #(1, 1'b0, 0, 0) c39148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39148));
	wire w118149;
	torch #(1'b1) c118149 (.i_clk(tick), .i_in(), .o_out(w118149));
	wire w134149;
	torch #(1'b1) c134149 (.i_clk(tick), .i_in(), .o_out(w134149));
	wire w152149;
	torch #(1'b1) c152149 (.i_clk(tick), .i_in(), .o_out(w152149));
	wire w168149;
	torch #(1'b1) c168149 (.i_clk(tick), .i_in(), .o_out(w168149));
	wire w125150;
	repeater #(2, 1'b0, 0, 0) c125150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125150));
	wire w159150;
	repeater #(2, 1'b0, 0, 0) c159150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159150));
	wire w48151;
	torch #(1'b1) c48151 (.i_clk(tick), .i_in(), .o_out(w48151));
	wire w52151;
	torch #(1'b1) c52151 (.i_clk(tick), .i_in(), .o_out(w52151));
	wire w56151;
	torch #(1'b1) c56151 (.i_clk(tick), .i_in(), .o_out(w56151));
	wire w60151;
	torch #(1'b1) c60151 (.i_clk(tick), .i_in(), .o_out(w60151));
	wire w119151;
	repeater #(2, 1'b0, 0, 0) c119151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119151));
	wire w135151;
	repeater #(1, 1'b0, 0, 0) c135151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135151));
	wire w153151;
	repeater #(2, 1'b0, 0, 0) c153151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153151));
	wire w169151;
	repeater #(1, 1'b0, 0, 0) c169151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169151));
	wire w129153;
	repeater #(1, 1'b0, 0, 0) c129153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w129153));
	wire w163153;
	repeater #(1, 1'b0, 0, 0) c163153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163153));
	wire w131154;
	repeater #(1, 1'b0, 0, 0) c131154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131154));
	wire w165154;
	repeater #(1, 1'b0, 0, 0) c165154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165154));
	wire w41155;
	torch #(1'b0) c41155 (.i_clk(tick), .i_in(), .o_out(w41155));
	wire w45155;
	torch #(1'b0) c45155 (.i_clk(tick), .i_in(), .o_out(w45155));
	wire w49155;
	torch #(1'b0) c49155 (.i_clk(tick), .i_in(), .o_out(w49155));
	wire w53155;
	torch #(1'b1) c53155 (.i_clk(tick), .i_in(), .o_out(w53155));
	wire w57155;
	torch #(1'b0) c57155 (.i_clk(tick), .i_in(), .o_out(w57155));
	wire w61155;
	torch #(1'b0) c61155 (.i_clk(tick), .i_in(), .o_out(w61155));
	wire w65155;
	torch #(1'b0) c65155 (.i_clk(tick), .i_in(), .o_out(w65155));
	wire w42157;
	torch #(1'b1) c42157 (.i_clk(tick), .i_in(), .o_out(w42157));
	wire w46157;
	torch #(1'b1) c46157 (.i_clk(tick), .i_in(), .o_out(w46157));
	wire w50157;
	torch #(1'b1) c50157 (.i_clk(tick), .i_in(), .o_out(w50157));
	wire w54157;
	torch #(1'b1) c54157 (.i_clk(tick), .i_in(), .o_out(w54157));
	wire w58157;
	torch #(1'b1) c58157 (.i_clk(tick), .i_in(), .o_out(w58157));
	wire w62157;
	torch #(1'b1) c62157 (.i_clk(tick), .i_in(), .o_out(w62157));
	wire w66157;
	torch #(1'b1) c66157 (.i_clk(tick), .i_in(), .o_out(w66157));
	wire w44162;

	wire w69162;
	repeater #(1, 1'b0, 0, 0) c69162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69162));
	wire w64163;

	wire w39164;
	repeater #(1, 1'b0, 0, 0) c39164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39164));
	wire w48167;
	torch #(1'b1) c48167 (.i_clk(tick), .i_in(), .o_out(w48167));
	wire w52167;
	torch #(1'b1) c52167 (.i_clk(tick), .i_in(), .o_out(w52167));
	wire w56167;
	torch #(1'b1) c56167 (.i_clk(tick), .i_in(), .o_out(w56167));
	wire w60167;
	torch #(1'b1) c60167 (.i_clk(tick), .i_in(), .o_out(w60167));
	wire w204167;

	wire w14168;

	wire w41171;
	torch #(1'b0) c41171 (.i_clk(tick), .i_in(), .o_out(w41171));
	wire w45171;
	torch #(1'b0) c45171 (.i_clk(tick), .i_in(), .o_out(w45171));
	wire w49171;
	torch #(1'b0) c49171 (.i_clk(tick), .i_in(), .o_out(w49171));
	wire w53171;
	torch #(1'b0) c53171 (.i_clk(tick), .i_in(), .o_out(w53171));
	wire w57171;
	torch #(1'b0) c57171 (.i_clk(tick), .i_in(), .o_out(w57171));
	wire w61171;
	torch #(1'b0) c61171 (.i_clk(tick), .i_in(), .o_out(w61171));
	wire w65171;
	torch #(1'b0) c65171 (.i_clk(tick), .i_in(), .o_out(w65171));
	wire w42173;
	torch #(1'b1) c42173 (.i_clk(tick), .i_in(), .o_out(w42173));
	wire w46173;
	torch #(1'b1) c46173 (.i_clk(tick), .i_in(), .o_out(w46173));
	wire w50173;
	torch #(1'b1) c50173 (.i_clk(tick), .i_in(), .o_out(w50173));
	wire w54173;
	torch #(1'b1) c54173 (.i_clk(tick), .i_in(), .o_out(w54173));
	wire w58173;
	torch #(1'b1) c58173 (.i_clk(tick), .i_in(), .o_out(w58173));
	wire w62173;
	torch #(1'b1) c62173 (.i_clk(tick), .i_in(), .o_out(w62173));
	wire w66173;
	torch #(1'b1) c66173 (.i_clk(tick), .i_in(), .o_out(w66173));
	wire w44178;

	wire w69178;
	repeater #(1, 1'b0, 0, 0) c69178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69178));
	wire w64179;

	wire w39180;
	repeater #(1, 1'b0, 0, 0) c39180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39180));
	wire w48183;
	torch #(1'b1) c48183 (.i_clk(tick), .i_in(), .o_out(w48183));
	wire w52183;
	torch #(1'b1) c52183 (.i_clk(tick), .i_in(), .o_out(w52183));
	wire w56183;
	torch #(1'b1) c56183 (.i_clk(tick), .i_in(), .o_out(w56183));
	wire w60183;
	torch #(1'b1) c60183 (.i_clk(tick), .i_in(), .o_out(w60183));
	wire w41187;
	torch #(1'b0) c41187 (.i_clk(tick), .i_in(), .o_out(w41187));
	wire w45187;
	torch #(1'b0) c45187 (.i_clk(tick), .i_in(), .o_out(w45187));
	wire w49187;
	torch #(1'b0) c49187 (.i_clk(tick), .i_in(), .o_out(w49187));
	wire w53187;
	torch #(1'b1) c53187 (.i_clk(tick), .i_in(), .o_out(w53187));
	wire w57187;
	torch #(1'b0) c57187 (.i_clk(tick), .i_in(), .o_out(w57187));
	wire w61187;
	torch #(1'b0) c61187 (.i_clk(tick), .i_in(), .o_out(w61187));
	wire w65187;
	torch #(1'b0) c65187 (.i_clk(tick), .i_in(), .o_out(w65187));
	wire w42189;
	torch #(1'b1) c42189 (.i_clk(tick), .i_in(), .o_out(w42189));
	wire w46189;
	torch #(1'b1) c46189 (.i_clk(tick), .i_in(), .o_out(w46189));
	wire w50189;
	torch #(1'b1) c50189 (.i_clk(tick), .i_in(), .o_out(w50189));
	wire w54189;
	torch #(1'b1) c54189 (.i_clk(tick), .i_in(), .o_out(w54189));
	wire w58189;
	torch #(1'b1) c58189 (.i_clk(tick), .i_in(), .o_out(w58189));
	wire w62189;
	torch #(1'b1) c62189 (.i_clk(tick), .i_in(), .o_out(w62189));
	wire w66189;
	torch #(1'b1) c66189 (.i_clk(tick), .i_in(), .o_out(w66189));
	wire w391101;
	repeater #(2, 1'b0, 0, 0) c391101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w391101));
	wire w431101;
	repeater #(2, 1'b0, 0, 0) c431101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w431101));
	wire w471101;
	repeater #(2, 1'b0, 0, 0) c471101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w471101));
	wire w511101;
	repeater #(2, 1'b0, 0, 0) c511101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w511101));
	wire w551101;
	repeater #(2, 1'b0, 0, 0) c551101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w551101));
	wire w591101;
	repeater #(2, 1'b0, 0, 0) c591101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w591101));
	wire w631101;
	repeater #(2, 1'b0, 0, 0) c631101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w631101));
	wire w401103;

	wire w441103;

	wire w481103;

	wire w521103;

	wire w561103;

	wire w601103;

	wire w641103;

	wire w401104;

	wire w441104;

	wire w481104;

	wire w521104;

	wire w561104;

	wire w601104;

	wire w641104;

	wire w391107;
	repeater #(1, 1'b1, 0, 0) c391107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w391107));
	wire w431107;
	repeater #(1, 1'b1, 0, 0) c431107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w431107));
	wire w471107;
	repeater #(1, 1'b1, 0, 0) c471107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w471107));
	wire w511107;
	repeater #(1, 1'b0, 0, 0) c511107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w511107));
	wire w551107;
	repeater #(1, 1'b1, 0, 0) c551107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w551107));
	wire w591107;
	repeater #(1, 1'b1, 0, 0) c591107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w591107));
	wire w631107;
	repeater #(1, 1'b1, 0, 0) c631107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w631107));
	wire w411108;

	wire w451108;

	wire w491108;

	wire w531108;

	wire w571108;

	wire w611108;

	wire w651108;

	wire w401109;

	wire w441109;

	wire w481109;

	wire w521109;

	wire w561109;

	wire w601109;

	wire w641109;

	wire w421111;
	torch #(1'b0) c421111 (.i_clk(tick), .i_in(), .o_out(w421111));
	wire w461111;
	torch #(1'b0) c461111 (.i_clk(tick), .i_in(), .o_out(w461111));
	wire w501111;
	torch #(1'b0) c501111 (.i_clk(tick), .i_in(), .o_out(w501111));
	wire w541111;
	torch #(1'b1) c541111 (.i_clk(tick), .i_in(), .o_out(w541111));
	wire w581111;
	torch #(1'b0) c581111 (.i_clk(tick), .i_in(), .o_out(w581111));
	wire w621111;
	torch #(1'b0) c621111 (.i_clk(tick), .i_in(), .o_out(w621111));
	wire w661111;
	torch #(1'b0) c661111 (.i_clk(tick), .i_in(), .o_out(w661111));
	wire w731124;
	repeater #(1, 1'b0, 0, 0) c731124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w731124));
	wire w122013;

	wire w155013;

	wire w156013;

	wire w189013;

	wire w190013;

	wire w15014;

	wire w16014;

	wire w49014;

	wire w123014;
	repeater #(1, 1'b1, 0, 0) c123014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123014));
	wire w157014;
	repeater #(1, 1'b1, 0, 0) c157014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157014));
	wire w191014;
	repeater #(1, 1'b1, 0, 0) c191014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191014));
	wire w17015;
	repeater #(1, 1'b1, 0, 0) c17015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17015));
	wire w120015;

	wire w153015;

	wire w154015;

	wire w187015;

	wire w188015;

	wire w13016;

	wire w14016;

	wire w47016;

	wire w50016;
	repeater #(1, 1'b1, 0, 0) c50016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50016));
	wire w121016;
	repeater #(1, 1'b1, 0, 0) c121016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121016));
	wire w155016;
	repeater #(1, 1'b1, 0, 0) c155016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155016));
	wire w189016;
	repeater #(1, 1'b1, 0, 0) c189016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189016));
	wire w15017;
	repeater #(1, 1'b1, 0, 0) c15017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15017));
	wire w49017;

	wire w118017;

	wire w151017;

	wire w152017;

	wire w185017;

	wire w186017;

	wire w11018;

	wire w12018;

	wire w45018;

	wire w48018;
	repeater #(1, 1'b1, 0, 0) c48018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48018));
	wire w119018;
	repeater #(1, 1'b1, 0, 0) c119018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119018));
	wire w153018;
	repeater #(1, 1'b1, 0, 0) c153018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153018));
	wire w187018;
	repeater #(1, 1'b1, 0, 0) c187018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187018));
	wire w13019;
	repeater #(1, 1'b1, 0, 0) c13019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13019));
	wire w47019;

	wire w116019;

	wire w149019;

	wire w150019;

	wire w183019;

	wire w184019;

	wire w9020;

	wire w10020;

	wire w43020;

	wire w46020;
	repeater #(1, 1'b1, 0, 0) c46020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46020));
	wire w117020;
	repeater #(1, 1'b1, 0, 0) c117020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117020));
	wire w151020;
	repeater #(1, 1'b1, 0, 0) c151020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151020));
	wire w185020;
	repeater #(1, 1'b1, 0, 0) c185020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185020));
	wire w11021;
	repeater #(1, 1'b1, 0, 0) c11021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11021));
	wire w45021;

	wire w114021;

	wire w147021;

	wire w148021;

	wire w181021;

	wire w182021;

	wire w7022;

	wire w8022;

	wire w41022;

	wire w44022;
	repeater #(1, 1'b1, 0, 0) c44022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44022));
	wire w115022;
	repeater #(1, 1'b1, 0, 0) c115022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115022));
	wire w149022;
	repeater #(1, 1'b1, 0, 0) c149022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149022));
	wire w183022;
	repeater #(1, 1'b1, 0, 0) c183022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183022));
	wire w9023;
	repeater #(1, 1'b1, 0, 0) c9023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9023));
	wire w43023;

	wire w112023;

	wire w145023;

	wire w146023;

	wire w179023;

	wire w180023;

	wire w5024;

	wire w6024;

	wire w39024;

	wire w42024;
	repeater #(1, 1'b1, 0, 0) c42024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42024));
	wire w113024;
	repeater #(1, 1'b1, 0, 0) c113024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113024));
	wire w147024;
	repeater #(1, 1'b1, 0, 0) c147024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147024));
	wire w181024;
	repeater #(1, 1'b1, 0, 0) c181024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181024));
	wire w7025;
	repeater #(1, 1'b1, 0, 0) c7025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7025));
	wire w41025;

	wire w110025;

	wire w143025;

	wire w144025;

	wire w177025;

	wire w178025;

	wire w3026;

	wire w4026;

	wire w37026;

	wire w40026;
	repeater #(1, 1'b1, 0, 0) c40026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40026));
	wire w111026;
	repeater #(1, 1'b1, 0, 0) c111026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111026));
	wire w145026;
	repeater #(1, 1'b1, 0, 0) c145026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145026));
	wire w179026;
	repeater #(1, 1'b1, 0, 0) c179026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179026));
	wire w5027;
	repeater #(1, 1'b1, 0, 0) c5027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5027));
	wire w39027;

	wire w108027;

	wire w141027;

	wire w142027;

	wire w175027;

	wire w176027;

	wire w1028;

	wire w2028;

	wire w35028;

	wire w38028;
	repeater #(1, 1'b1, 0, 0) c38028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38028));
	wire w109028;
	repeater #(1, 1'b0, 0, 0) c109028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109028));
	wire w143028;
	repeater #(1, 1'b0, 0, 0) c143028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143028));
	wire w177028;
	repeater #(1, 1'b0, 0, 0) c177028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177028));
	wire w3029;
	repeater #(1, 1'b0, 0, 0) c3029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3029));
	wire w37029;

	wire w106029;

	wire w139029;

	wire w140029;

	wire w173029;

	wire w174029;

	wire w207029;

	wire w0030;

	wire w33030;

	wire w36030;
	repeater #(1, 1'b0, 0, 0) c36030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36030));
	wire w107030;
	repeater #(1, 1'b1, 0, 0) c107030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107030));
	wire w141030;
	repeater #(1, 1'b1, 0, 0) c141030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141030));
	wire w175030;
	repeater #(1, 1'b1, 0, 0) c175030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175030));
	wire w1031;
	repeater #(1, 1'b1, 0, 0) c1031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1031));
	wire w35031;

	wire w104031;

	wire w137031;

	wire w138031;

	wire w171031;

	wire w172031;

	wire w205031;

	wire w206031;

	wire w31032;

	wire w34032;
	repeater #(1, 1'b1, 0, 0) c34032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34032));
	wire w105032;
	repeater #(1, 1'b1, 0, 0) c105032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105032));
	wire w139032;
	repeater #(1, 1'b1, 0, 0) c139032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139032));
	wire w173032;
	repeater #(1, 1'b1, 0, 0) c173032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173032));
	wire w207032;
	repeater #(1, 1'b1, 0, 0) c207032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207032));
	wire w33033;

	wire w102033;

	wire w135033;

	wire w136033;

	wire w169033;

	wire w170033;

	wire w203033;

	wire w204033;

	wire w29034;

	wire w32034;
	repeater #(1, 1'b1, 0, 0) c32034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32034));
	wire w103034;
	repeater #(1, 1'b1, 0, 0) c103034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103034));
	wire w137034;
	repeater #(1, 1'b1, 0, 0) c137034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137034));
	wire w171034;
	repeater #(1, 1'b1, 0, 0) c171034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171034));
	wire w205034;
	repeater #(1, 1'b1, 0, 0) c205034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205034));
	wire w31035;

	wire w100035;

	wire w133035;

	wire w134035;

	wire w167035;

	wire w168035;

	wire w201035;

	wire w202035;

	wire w27036;

	wire w30036;
	repeater #(1, 1'b1, 0, 0) c30036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30036));
	wire w101036;
	repeater #(1, 1'b1, 0, 0) c101036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101036));
	wire w135036;
	repeater #(1, 1'b1, 0, 0) c135036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135036));
	wire w169036;
	repeater #(1, 1'b1, 0, 0) c169036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169036));
	wire w203036;
	repeater #(1, 1'b1, 0, 0) c203036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203036));
	wire w29037;

	wire w98037;

	wire w131037;

	wire w132037;

	wire w165037;

	wire w166037;

	wire w199037;

	wire w200037;

	wire w25038;

	wire w28038;
	repeater #(1, 1'b1, 0, 0) c28038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28038));
	wire w99038;
	repeater #(1, 1'b1, 0, 0) c99038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99038));
	wire w133038;
	repeater #(1, 1'b1, 0, 0) c133038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133038));
	wire w167038;
	repeater #(1, 1'b1, 0, 0) c167038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167038));
	wire w201038;
	repeater #(1, 1'b1, 0, 0) c201038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201038));
	wire w27039;

	wire w129039;

	wire w163039;

	wire w197039;

	wire w23040;

	wire w26040;
	repeater #(1, 1'b1, 0, 0) c26040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26040));
	wire w97040;
	repeater #(1, 1'b1, 0, 0) c97040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97040));
	wire w131040;
	repeater #(1, 1'b1, 0, 0) c131040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131040));
	wire w165040;
	repeater #(1, 1'b1, 0, 0) c165040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165040));
	wire w199040;
	repeater #(1, 1'b1, 0, 0) c199040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199040));
	wire w25041;

	wire w24042;
	repeater #(2, 1'b1, 0, 0) c24042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24042));
	wire w26043;
	repeater #(1, 1'b1, 0, 0) c26043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26043));
	wire w116045;
	repeater #(2, 1'b1, 0, 0) c116045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116045));
	wire w150045;
	repeater #(2, 1'b1, 0, 0) c150045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150045));
	wire w25046;
	torch #(1'b1) c25046 (.i_clk(tick), .i_in(), .o_out(w25046));
	wire w29046;
	torch #(1'b1) c29046 (.i_clk(tick), .i_in(), .o_out(w29046));
	wire w33046;
	torch #(1'b1) c33046 (.i_clk(tick), .i_in(), .o_out(w33046));
	wire w37046;
	torch #(1'b0) c37046 (.i_clk(tick), .i_in(), .o_out(w37046));
	wire w41046;
	torch #(1'b1) c41046 (.i_clk(tick), .i_in(), .o_out(w41046));
	wire w45046;
	torch #(1'b1) c45046 (.i_clk(tick), .i_in(), .o_out(w45046));
	wire w49046;
	torch #(1'b1) c49046 (.i_clk(tick), .i_in(), .o_out(w49046));
	wire w102047;
	repeater #(1, 1'b1, 0, 0) c102047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102047));
	wire w108047;
	torch #(1'b1) c108047 (.i_clk(tick), .i_in(), .o_out(w108047));
	wire w118047;
	repeater #(1, 1'b1, 0, 0) c118047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118047));
	wire w136047;
	repeater #(1, 1'b1, 0, 0) c136047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136047));
	wire w142047;
	torch #(1'b1) c142047 (.i_clk(tick), .i_in(), .o_out(w142047));
	wire w152047;
	repeater #(1, 1'b1, 0, 0) c152047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152047));
	wire w26049;
	repeater #(1, 1'b1, 0, 0) c26049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26049));
	wire w30049;
	repeater #(1, 1'b1, 0, 0) c30049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30049));
	wire w34049;
	repeater #(1, 1'b1, 0, 0) c34049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34049));
	wire w38049;
	repeater #(1, 1'b0, 0, 0) c38049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38049));
	wire w42049;
	repeater #(1, 1'b1, 0, 0) c42049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42049));
	wire w46049;
	repeater #(1, 1'b1, 0, 0) c46049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46049));
	wire w50049;
	repeater #(1, 1'b1, 0, 0) c50049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50049));
	wire w25050;
	torch #(1'b1) c25050 (.i_clk(tick), .i_in(), .o_out(w25050));
	wire w29050;
	torch #(1'b1) c29050 (.i_clk(tick), .i_in(), .o_out(w29050));
	wire w33050;
	torch #(1'b1) c33050 (.i_clk(tick), .i_in(), .o_out(w33050));
	wire w37050;
	torch #(1'b0) c37050 (.i_clk(tick), .i_in(), .o_out(w37050));
	wire w41050;
	torch #(1'b1) c41050 (.i_clk(tick), .i_in(), .o_out(w41050));
	wire w45050;
	torch #(1'b1) c45050 (.i_clk(tick), .i_in(), .o_out(w45050));
	wire w49050;
	torch #(1'b1) c49050 (.i_clk(tick), .i_in(), .o_out(w49050));
	wire w109050;
	repeater #(1, 1'b1, 0, 0) c109050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109050));
	wire w143050;
	repeater #(1, 1'b1, 0, 0) c143050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143050));
	wire w102051;
	repeater #(1, 1'b1, 0, 0) c102051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102051));
	wire w118051;
	repeater #(1, 1'b1, 0, 0) c118051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118051));
	wire w136051;
	repeater #(1, 1'b1, 0, 0) c136051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136051));
	wire w152051;
	repeater #(1, 1'b1, 0, 0) c152051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152051));
	wire w171051;
	torch #(1'b1) c171051 (.i_clk(tick), .i_in(), .o_out(w171051));
	wire w175051;
	torch #(1'b1) c175051 (.i_clk(tick), .i_in(), .o_out(w175051));
	wire w179051;
	torch #(1'b0) c179051 (.i_clk(tick), .i_in(), .o_out(w179051));
	wire w183051;
	torch #(1'b0) c183051 (.i_clk(tick), .i_in(), .o_out(w183051));
	wire w207051;
	torch #(1'b0) c207051 (.i_clk(tick), .i_in(), .o_out(w207051));
	wire w3052;
	torch #(1'b0) c3052 (.i_clk(tick), .i_in(), .o_out(w3052));
	wire w7052;
	torch #(1'b0) c7052 (.i_clk(tick), .i_in(), .o_out(w7052));
	wire w11052;
	torch #(1'b0) c11052 (.i_clk(tick), .i_in(), .o_out(w11052));
	wire w107052;

	wire w141052;

	wire w24053;
	torch #(1'b0) c24053 (.i_clk(tick), .i_in(), .o_out(w24053));
	wire w28053;
	torch #(1'b0) c28053 (.i_clk(tick), .i_in(), .o_out(w28053));
	wire w32053;
	torch #(1'b0) c32053 (.i_clk(tick), .i_in(), .o_out(w32053));
	wire w36053;
	torch #(1'b1) c36053 (.i_clk(tick), .i_in(), .o_out(w36053));
	wire w40053;
	torch #(1'b0) c40053 (.i_clk(tick), .i_in(), .o_out(w40053));
	wire w44053;
	torch #(1'b0) c44053 (.i_clk(tick), .i_in(), .o_out(w44053));
	wire w48053;
	torch #(1'b0) c48053 (.i_clk(tick), .i_in(), .o_out(w48053));
	wire w115053;

	wire w149053;

	wire w101054;

	wire w102054;

	wire w112054;

	wire w117054;

	wire w118054;

	wire w135054;

	wire w136054;

	wire w146054;

	wire w151054;

	wire w152054;

	wire w94056;

	wire w110056;

	wire w128056;

	wire w144056;

	wire w100057;

	wire w101057;

	wire w116057;

	wire w117057;

	wire w134057;

	wire w135057;

	wire w150057;

	wire w151057;

	wire w110058;

	wire w144058;

	wire w173058;
	repeater #(1, 1'b1, 0, 0) c173058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173058));
	wire w175058;
	repeater #(2, 1'b0, 0, 0) c175058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175058));
	wire w177058;
	repeater #(2, 1'b0, 0, 0) c177058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177058));
	wire w181058;
	repeater #(2, 1'b1, 0, 0) c181058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181058));
	wire w183058;
	repeater #(2, 1'b1, 0, 0) c183058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183058));
	wire w185058;
	repeater #(1, 1'b1, 0, 0) c185058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185058));
	wire w205058;
	repeater #(1, 1'b1, 0, 0) c205058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205058));
	wire w207058;
	repeater #(2, 1'b1, 0, 0) c207058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207058));
	wire w1059;
	repeater #(2, 1'b1, 0, 0) c1059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1059));
	wire w5059;
	repeater #(2, 1'b1, 0, 0) c5059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5059));
	wire w7059;
	repeater #(2, 1'b1, 0, 0) c7059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7059));
	wire w9059;
	repeater #(1, 1'b1, 0, 0) c9059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9059));
	wire w32059;
	torch #(1'b1) c32059 (.i_clk(tick), .i_in(), .o_out(w32059));
	wire w36059;
	torch #(1'b1) c36059 (.i_clk(tick), .i_in(), .o_out(w36059));
	wire w40059;
	torch #(1'b1) c40059 (.i_clk(tick), .i_in(), .o_out(w40059));
	wire w44059;
	torch #(1'b1) c44059 (.i_clk(tick), .i_in(), .o_out(w44059));
	wire w170059;
	repeater #(1, 1'b1, 0, 0) c170059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170059));
	wire w12060;
	repeater #(1, 1'b1, 0, 0) c12060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12060));
	wire w53060;
	repeater #(1, 1'b0, 0, 0) c53060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53060));
	wire w94060;

	wire w98060;

	wire w102060;

	wire w106060;

	wire w110060;

	wire w114060;

	wire w118060;

	wire w128060;

	wire w132060;

	wire w136060;

	wire w140060;

	wire w144060;

	wire w148060;

	wire w152060;

	wire w180060;

	wire w2061;

	wire w172061;

	wire w176061;

	wire w179061;

	wire w181061;

	wire w184061;

	wire w206061;

	wire w1062;

	wire w3062;

	wire w6062;

	wire w10062;

	wire w171062;

	wire w173062;

	wire w175062;

	wire w177062;

	wire w180062;

	wire w183062;

	wire w185062;

	wire w205062;

	wire w207062;

	wire w2063;

	wire w5063;

	wire w7063;

	wire w9063;

	wire w11063;

	wire w176063;

	wire w6064;

	wire w94064;

	wire w98064;

	wire w102064;

	wire w106064;

	wire w110064;

	wire w114064;

	wire w118064;

	wire w128064;

	wire w132064;

	wire w136064;

	wire w140064;

	wire w144064;

	wire w148064;

	wire w152064;

	wire w172064;

	wire w176064;

	wire w177064;

	wire w181064;

	wire w183064;

	wire w185064;

	wire w205064;

	wire w207064;

	wire w1065;

	wire w5065;

	wire w6065;

	wire w10065;

	wire w177065;

	wire w5066;

	wire w92066;
	repeater #(1, 1'b1, 0, 0) c92066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92066));
	wire w96066;
	repeater #(1, 1'b1, 0, 0) c96066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96066));
	wire w100066;
	repeater #(1, 1'b1, 0, 0) c100066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100066));
	wire w104066;
	repeater #(1, 1'b1, 0, 0) c104066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104066));
	wire w126066;
	repeater #(1, 1'b1, 0, 0) c126066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126066));
	wire w130066;
	repeater #(1, 1'b1, 0, 0) c130066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130066));
	wire w134066;
	repeater #(1, 1'b1, 0, 0) c134066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134066));
	wire w138066;
	repeater #(1, 1'b1, 0, 0) c138066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138066));
	wire w167066;
	repeater #(1, 1'b1, 0, 0) c167066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167066));
	wire w172066;
	repeater #(1, 1'b1, 0, 0) c172066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172066));
	wire w175066;
	repeater #(2, 1'b1, 0, 0) c175066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175066));
	wire w177066;

	wire w5067;

	wire w7067;
	repeater #(2, 1'b1, 0, 0) c7067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7067));
	wire w10067;
	repeater #(1, 1'b1, 0, 0) c10067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10067));
	wire w15067;
	repeater #(1, 1'b1, 0, 0) c15067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15067));
	wire w110067;

	wire w114067;

	wire w118067;

	wire w144067;

	wire w148067;

	wire w152067;

	wire w166067;

	wire w167067;
	repeater #(1, 1'b1, 0, 0) c167067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167067));
	wire w171067;

	wire w172067;
	repeater #(1, 1'b1, 0, 0) c172067 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172067));
	wire w178067;

	wire w4068;

	wire w10068;
	repeater #(1, 1'b1, 0, 0) c10068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10068));
	wire w11068;

	wire w15068;
	repeater #(1, 1'b1, 0, 0) c15068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15068));
	wire w16068;

	wire w25068;
	torch #(1'b1) c25068 (.i_clk(tick), .i_in(), .o_out(w25068));
	wire w29068;
	torch #(1'b1) c29068 (.i_clk(tick), .i_in(), .o_out(w29068));
	wire w33068;
	torch #(1'b1) c33068 (.i_clk(tick), .i_in(), .o_out(w33068));
	wire w37068;
	torch #(1'b0) c37068 (.i_clk(tick), .i_in(), .o_out(w37068));
	wire w41068;
	torch #(1'b1) c41068 (.i_clk(tick), .i_in(), .o_out(w41068));
	wire w45068;
	torch #(1'b1) c45068 (.i_clk(tick), .i_in(), .o_out(w45068));
	wire w49068;
	torch #(1'b1) c49068 (.i_clk(tick), .i_in(), .o_out(w49068));
	wire w26069;
	repeater #(1, 1'b0, 0, 0) c26069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26069));
	wire w30069;
	repeater #(1, 1'b0, 0, 0) c30069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30069));
	wire w34069;
	repeater #(1, 1'b0, 0, 0) c34069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34069));
	wire w38069;
	repeater #(1, 1'b1, 0, 0) c38069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38069));
	wire w42069;
	repeater #(1, 1'b0, 0, 0) c42069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42069));
	wire w46069;
	repeater #(1, 1'b0, 0, 0) c46069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46069));
	wire w50069;
	repeater #(1, 1'b0, 0, 0) c50069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50069));
	wire w110069;

	wire w144069;

	wire w92070;
	repeater #(1, 1'b1, 0, 0) c92070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92070));
	wire w108070;
	repeater #(1, 1'b1, 0, 0) c108070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108070));
	wire w126070;
	repeater #(1, 1'b1, 0, 0) c126070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126070));
	wire w142070;
	repeater #(1, 1'b1, 0, 0) c142070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142070));
	wire w167070;
	repeater #(1, 1'b1, 0, 0) c167070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167070));
	wire w172070;
	repeater #(1, 1'b1, 0, 0) c172070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172070));
	wire w177070;
	repeater #(1, 1'b1, 0, 0) c177070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177070));
	wire w5071;
	repeater #(1, 1'b1, 0, 0) c5071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5071));
	wire w10071;
	repeater #(1, 1'b1, 0, 0) c10071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10071));
	wire w15071;
	repeater #(1, 1'b1, 0, 0) c15071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15071));
	wire w24071;

	wire w26071;
	repeater #(1, 1'b0, 0, 0) c26071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26071));
	wire w28071;

	wire w30071;
	repeater #(1, 1'b0, 0, 0) c30071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30071));
	wire w32071;

	wire w34071;
	repeater #(1, 1'b0, 0, 0) c34071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34071));
	wire w36071;

	wire w38071;
	repeater #(1, 1'b1, 0, 0) c38071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38071));
	wire w40071;

	wire w42071;
	repeater #(1, 1'b0, 0, 0) c42071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42071));
	wire w44071;

	wire w46071;
	repeater #(1, 1'b0, 0, 0) c46071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46071));
	wire w48071;

	wire w50071;
	repeater #(1, 1'b0, 0, 0) c50071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50071));
	wire w99071;
	repeater #(1, 1'b1, 0, 0) c99071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99071));
	wire w115071;
	repeater #(1, 1'b1, 0, 0) c115071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115071));
	wire w133071;
	repeater #(1, 1'b1, 0, 0) c133071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133071));
	wire w149071;
	repeater #(1, 1'b1, 0, 0) c149071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149071));
	wire w166071;

	wire w167071;
	repeater #(1, 1'b1, 0, 0) c167071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167071));
	wire w171071;

	wire w172071;
	repeater #(1, 1'b1, 0, 0) c172071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172071));
	wire w176071;

	wire w177071;
	repeater #(1, 1'b1, 0, 0) c177071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177071));
	wire w5072;
	repeater #(1, 1'b1, 0, 0) c5072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5072));
	wire w6072;

	wire w10072;
	repeater #(1, 1'b1, 0, 0) c10072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10072));
	wire w11072;

	wire w15072;
	repeater #(1, 1'b1, 0, 0) c15072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15072));
	wire w16072;

	wire w94072;

	wire w110072;

	wire w128072;

	wire w144072;

	wire w102073;

	wire w136073;

	wire w97074;

	wire w99074;

	wire w100074;

	wire w105074;

	wire w113074;

	wire w115074;

	wire w131074;

	wire w133074;

	wire w134074;

	wire w139074;

	wire w147074;

	wire w149074;

	wire w167074;
	repeater #(1, 1'b0, 0, 0) c167074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167074));
	wire w172074;
	repeater #(1, 1'b0, 0, 0) c172074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172074));
	wire w177074;
	repeater #(1, 1'b1, 0, 0) c177074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177074));
	wire w5075;
	repeater #(1, 1'b1, 0, 0) c5075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5075));
	wire w10075;
	repeater #(1, 1'b0, 0, 0) c10075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10075));
	wire w15075;
	repeater #(1, 1'b0, 0, 0) c15075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15075));
	wire w32075;
	torch #(1'b1) c32075 (.i_clk(tick), .i_in(), .o_out(w32075));
	wire w36075;
	torch #(1'b1) c36075 (.i_clk(tick), .i_in(), .o_out(w36075));
	wire w40075;
	torch #(1'b1) c40075 (.i_clk(tick), .i_in(), .o_out(w40075));
	wire w44075;
	torch #(1'b1) c44075 (.i_clk(tick), .i_in(), .o_out(w44075));
	wire w166075;

	wire w167075;
	repeater #(1, 1'b0, 0, 0) c167075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167075));
	wire w171075;

	wire w172075;
	repeater #(1, 1'b0, 0, 0) c172075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172075));
	wire w176075;

	wire w177075;
	repeater #(1, 1'b1, 0, 0) c177075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177075));
	wire w5076;
	repeater #(1, 1'b1, 0, 0) c5076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5076));
	wire w6076;

	wire w10076;
	repeater #(1, 1'b0, 0, 0) c10076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10076));
	wire w11076;

	wire w15076;
	repeater #(1, 1'b0, 0, 0) c15076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15076));
	wire w16076;

	wire w53076;
	repeater #(1, 1'b0, 0, 0) c53076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53076));
	wire w107076;

	wire w108076;

	wire w141076;

	wire w142076;

	wire w97078;

	wire w99078;

	wire w100078;

	wire w113078;

	wire w115078;

	wire w116078;

	wire w131078;

	wire w133078;

	wire w134078;

	wire w147078;

	wire w149078;

	wire w150078;

	wire w167078;
	repeater #(1, 1'b0, 0, 0) c167078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167078));
	wire w172078;
	repeater #(1, 1'b0, 0, 0) c172078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172078));
	wire w177078;
	repeater #(1, 1'b0, 0, 0) c177078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177078));
	wire w5079;
	repeater #(1, 1'b0, 0, 0) c5079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5079));
	wire w10079;
	repeater #(1, 1'b0, 0, 0) c10079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10079));
	wire w15079;
	repeater #(1, 1'b0, 0, 0) c15079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15079));
	wire w166079;

	wire w167079;
	repeater #(1, 1'b0, 0, 0) c167079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167079));
	wire w171079;

	wire w172079;
	repeater #(1, 1'b0, 0, 0) c172079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172079));
	wire w176079;

	wire w177079;
	repeater #(1, 1'b0, 0, 0) c177079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177079));
	wire w184079;
	repeater #(1, 1'b0, 0, 0) c184079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184079));
	wire w206079;
	repeater #(1, 1'b0, 0, 0) c206079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206079));
	wire w5080;
	repeater #(1, 1'b0, 0, 0) c5080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5080));
	wire w6080;

	wire w10080;
	repeater #(1, 1'b0, 0, 0) c10080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10080));
	wire w11080;

	wire w15080;
	repeater #(1, 1'b0, 0, 0) c15080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15080));
	wire w16080;

	wire w94080;
	torch #(1'b1) c94080 (.i_clk(tick), .i_in(), .o_out(w94080));
	wire w95080;

	wire w110080;
	torch #(1'b1) c110080 (.i_clk(tick), .i_in(), .o_out(w110080));
	wire w111080;

	wire w128080;
	torch #(1'b1) c128080 (.i_clk(tick), .i_in(), .o_out(w128080));
	wire w129080;

	wire w144080;
	torch #(1'b1) c144080 (.i_clk(tick), .i_in(), .o_out(w144080));
	wire w145080;

	wire w168080;
	repeater #(2, 1'b1, 0, 0) c168080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168080));
	wire w177080;
	repeater #(2, 1'b0, 0, 0) c177080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177080));
	wire w195080;

	wire w5081;
	repeater #(2, 1'b0, 0, 0) c5081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5081));
	wire w14081;
	repeater #(2, 1'b1, 0, 0) c14081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14081));
	wire w95081;

	wire w97081;

	wire w111081;

	wire w113081;

	wire w129081;

	wire w131081;

	wire w145081;

	wire w147081;

	wire w166081;

	wire w167081;

	wire w173081;
	repeater #(1, 1'b0, 0, 0) c173081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173081));
	wire w174081;
	repeater #(2, 1'b0, 0, 0) c174081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174081));
	wire w196081;

	wire w8082;
	repeater #(2, 1'b0, 0, 0) c8082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8082));
	wire w9082;
	repeater #(1, 1'b0, 0, 0) c9082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9082));
	wire w15082;

	wire w16082;

	wire w170082;
	repeater #(2, 1'b0, 0, 0) c170082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170082));
	wire w171082;
	repeater #(2, 1'b0, 0, 0) c171082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171082));
	wire w173082;

	wire w187082;
	repeater #(1, 1'b1, 0, 0) c187082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187082));
	wire w188082;

	wire w196082;
	repeater #(1, 1'b0, 0, 0) c196082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196082));
	wire w202082;

	wire w203082;
	repeater #(1, 1'b1, 0, 0) c203082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203082));
	wire w9083;

	wire w11083;
	repeater #(2, 1'b0, 0, 0) c11083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11083));
	wire w12083;
	repeater #(2, 1'b0, 0, 0) c12083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12083));
	wire w97083;

	wire w98083;

	wire w99083;

	wire w113083;

	wire w114083;

	wire w115083;

	wire w131083;

	wire w132083;

	wire w133083;

	wire w147083;

	wire w148083;

	wire w149083;

	wire w171083;

	wire w173083;
	repeater #(1, 1'b0, 0, 0) c173083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173083));
	wire w184083;

	wire w185083;

	wire w205083;

	wire w206083;

	wire w9084;
	repeater #(1, 1'b1, 0, 0) c9084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9084));
	wire w11084;

	wire w25084;
	torch #(1'b1) c25084 (.i_clk(tick), .i_in(), .o_out(w25084));
	wire w29084;
	torch #(1'b1) c29084 (.i_clk(tick), .i_in(), .o_out(w29084));
	wire w33084;
	torch #(1'b1) c33084 (.i_clk(tick), .i_in(), .o_out(w33084));
	wire w37084;
	torch #(1'b1) c37084 (.i_clk(tick), .i_in(), .o_out(w37084));
	wire w41084;
	torch #(1'b1) c41084 (.i_clk(tick), .i_in(), .o_out(w41084));
	wire w45084;
	torch #(1'b1) c45084 (.i_clk(tick), .i_in(), .o_out(w45084));
	wire w49084;
	torch #(1'b1) c49084 (.i_clk(tick), .i_in(), .o_out(w49084));
	wire w99084;

	wire w108084;

	wire w109084;

	wire w115084;

	wire w133084;

	wire w142084;

	wire w143084;

	wire w149084;

	wire w167084;

	wire w171084;

	wire w195084;

	wire w196084;

	wire w11085;

	wire w15085;

	wire w26085;
	repeater #(1, 1'b0, 0, 0) c26085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26085));
	wire w30085;
	repeater #(1, 1'b0, 0, 0) c30085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30085));
	wire w34085;
	repeater #(1, 1'b0, 0, 0) c34085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34085));
	wire w38085;
	repeater #(1, 1'b1, 0, 0) c38085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38085));
	wire w42085;
	repeater #(1, 1'b0, 0, 0) c42085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42085));
	wire w46085;
	repeater #(1, 1'b0, 0, 0) c46085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46085));
	wire w50085;
	repeater #(1, 1'b0, 0, 0) c50085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50085));
	wire w167085;

	wire w169085;
	repeater #(1, 1'b0, 0, 0) c169085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169085));
	wire w174085;

	wire w178085;

	wire w184085;
	repeater #(1, 1'b0, 0, 0) c184085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184085));
	wire w192085;

	wire w193085;
	repeater #(1, 1'b0, 0, 0) c193085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193085));
	wire w206085;
	repeater #(1, 1'b0, 0, 0) c206085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206085));
	wire w4086;

	wire w8086;

	wire w13086;
	repeater #(1, 1'b1, 0, 0) c13086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13086));
	wire w15086;

	wire w97086;
	repeater #(1, 1'b0, 0, 0) c97086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97086));
	wire w99086;
	torch #(1'b0) c99086 (.i_clk(tick), .i_in(), .o_out(w99086));
	wire w105086;
	torch #(1'b0) c105086 (.i_clk(tick), .i_in(), .o_out(w105086));
	wire w113086;
	repeater #(1, 1'b0, 0, 0) c113086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113086));
	wire w115086;
	torch #(1'b0) c115086 (.i_clk(tick), .i_in(), .o_out(w115086));
	wire w121086;
	torch #(1'b0) c121086 (.i_clk(tick), .i_in(), .o_out(w121086));
	wire w131086;
	repeater #(1, 1'b0, 0, 0) c131086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131086));
	wire w133086;
	torch #(1'b0) c133086 (.i_clk(tick), .i_in(), .o_out(w133086));
	wire w139086;
	torch #(1'b0) c139086 (.i_clk(tick), .i_in(), .o_out(w139086));
	wire w147086;
	repeater #(1, 1'b0, 0, 0) c147086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147086));
	wire w149086;
	torch #(1'b0) c149086 (.i_clk(tick), .i_in(), .o_out(w149086));
	wire w155086;
	torch #(1'b0) c155086 (.i_clk(tick), .i_in(), .o_out(w155086));
	wire w174086;

	wire w176086;
	repeater #(1, 1'b0, 0, 0) c176086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176086));
	wire w177086;

	wire w184086;

	wire w201086;

	wire w206086;

	wire w5087;

	wire w6087;
	repeater #(1, 1'b1, 0, 0) c6087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6087));
	wire w8087;

	wire w24087;

	wire w26087;
	repeater #(1, 1'b0, 0, 0) c26087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26087));
	wire w28087;

	wire w30087;
	repeater #(1, 1'b0, 0, 0) c30087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30087));
	wire w32087;

	wire w34087;
	repeater #(1, 1'b0, 0, 0) c34087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34087));
	wire w36087;

	wire w38087;
	repeater #(1, 1'b1, 0, 0) c38087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38087));
	wire w40087;

	wire w42087;
	repeater #(1, 1'b0, 0, 0) c42087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42087));
	wire w44087;

	wire w46087;
	repeater #(1, 1'b0, 0, 0) c46087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46087));
	wire w48087;

	wire w50087;
	repeater #(1, 1'b0, 0, 0) c50087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50087));
	wire w170087;

	wire w185087;

	wire w189087;
	repeater #(1, 1'b0, 0, 0) c189087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189087));
	wire w202087;
	repeater #(2, 1'b1, 0, 0) c202087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202087));
	wire w205087;

	wire w12088;

	wire w101088;
	repeater #(1, 1'b1, 0, 0) c101088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101088));
	wire w117088;
	repeater #(1, 1'b1, 0, 0) c117088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117088));
	wire w135088;
	repeater #(1, 1'b1, 0, 0) c135088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135088));
	wire w151088;
	repeater #(1, 1'b1, 0, 0) c151088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151088));
	wire w167088;

	wire w168088;
	repeater #(1, 1'b0, 0, 0) c168088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168088));
	wire w175088;
	repeater #(2, 1'b0, 0, 0) c175088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175088));
	wire w188088;
	assign outputs[56] = ();
	wire w7089;
	repeater #(2, 1'b1, 0, 0) c7089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7089));
	wire w14089;
	repeater #(1, 1'b0, 0, 0) c14089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14089));
	wire w15089;

	wire w98090;
	torch #(1'b1) c98090 (.i_clk(tick), .i_in(), .o_out(w98090));
	wire w114090;
	torch #(1'b1) c114090 (.i_clk(tick), .i_in(), .o_out(w114090));
	wire w132090;
	torch #(1'b1) c132090 (.i_clk(tick), .i_in(), .o_out(w132090));
	wire w148090;
	torch #(1'b1) c148090 (.i_clk(tick), .i_in(), .o_out(w148090));
	wire w32091;
	torch #(1'b1) c32091 (.i_clk(tick), .i_in(), .o_out(w32091));
	wire w36091;
	torch #(1'b1) c36091 (.i_clk(tick), .i_in(), .o_out(w36091));
	wire w40091;
	torch #(1'b1) c40091 (.i_clk(tick), .i_in(), .o_out(w40091));
	wire w44091;
	torch #(1'b1) c44091 (.i_clk(tick), .i_in(), .o_out(w44091));
	wire w53092;
	repeater #(1, 1'b0, 0, 0) c53092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53092));
	wire w106092;
	torch #(1'b1) c106092 (.i_clk(tick), .i_in(), .o_out(w106092));
	wire w122092;
	torch #(1'b1) c122092 (.i_clk(tick), .i_in(), .o_out(w122092));
	wire w140092;
	torch #(1'b1) c140092 (.i_clk(tick), .i_in(), .o_out(w140092));
	wire w156092;
	torch #(1'b1) c156092 (.i_clk(tick), .i_in(), .o_out(w156092));
	wire w97093;
	repeater #(2, 1'b0, 0, 0) c97093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97093));
	wire w113093;
	repeater #(2, 1'b0, 0, 0) c113093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113093));
	wire w131093;
	repeater #(2, 1'b0, 0, 0) c131093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131093));
	wire w147093;
	repeater #(2, 1'b0, 0, 0) c147093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147093));
	wire w107094;
	repeater #(2, 1'b0, 0, 0) c107094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107094));
	wire w123094;
	repeater #(1, 1'b0, 0, 0) c123094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123094));
	wire w141094;
	repeater #(2, 1'b0, 0, 0) c141094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141094));
	wire w157094;
	repeater #(1, 1'b0, 0, 0) c157094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157094));
	wire w117096;
	repeater #(1, 1'b0, 0, 0) c117096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117096));
	wire w151096;
	repeater #(1, 1'b0, 0, 0) c151096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151096));
	wire w119097;
	repeater #(1, 1'b0, 0, 0) c119097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119097));
	wire w153097;
	repeater #(1, 1'b0, 0, 0) c153097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153097));
	wire w250100;
	torch #(1'b1) c250100 (.i_clk(tick), .i_in(), .o_out(w250100));
	wire w290100;
	torch #(1'b1) c290100 (.i_clk(tick), .i_in(), .o_out(w290100));
	wire w330100;
	torch #(1'b1) c330100 (.i_clk(tick), .i_in(), .o_out(w330100));
	wire w370100;
	torch #(1'b0) c370100 (.i_clk(tick), .i_in(), .o_out(w370100));
	wire w410100;
	torch #(1'b1) c410100 (.i_clk(tick), .i_in(), .o_out(w410100));
	wire w450100;
	torch #(1'b1) c450100 (.i_clk(tick), .i_in(), .o_out(w450100));
	wire w490100;
	torch #(1'b1) c490100 (.i_clk(tick), .i_in(), .o_out(w490100));
	wire w260101;
	repeater #(1, 1'b0, 0, 0) c260101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260101));
	wire w300101;
	repeater #(1, 1'b0, 0, 0) c300101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300101));
	wire w340101;
	repeater #(1, 1'b0, 0, 0) c340101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340101));
	wire w380101;
	repeater #(1, 1'b1, 0, 0) c380101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380101));
	wire w420101;
	repeater #(1, 1'b0, 0, 0) c420101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420101));
	wire w460101;
	repeater #(1, 1'b0, 0, 0) c460101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460101));
	wire w500101;
	repeater #(1, 1'b0, 0, 0) c500101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500101));
	wire w240103;

	wire w260103;
	repeater #(1, 1'b0, 0, 0) c260103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260103));
	wire w280103;

	wire w300103;
	repeater #(1, 1'b0, 0, 0) c300103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300103));
	wire w320103;

	wire w340103;
	repeater #(1, 1'b0, 0, 0) c340103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340103));
	wire w360103;

	wire w380103;
	repeater #(1, 1'b1, 0, 0) c380103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380103));
	wire w400103;

	wire w420103;
	repeater #(1, 1'b0, 0, 0) c420103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420103));
	wire w440103;

	wire w460103;
	repeater #(1, 1'b0, 0, 0) c460103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460103));
	wire w480103;

	wire w500103;
	repeater #(1, 1'b0, 0, 0) c500103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500103));
	wire w320107;
	torch #(1'b1) c320107 (.i_clk(tick), .i_in(), .o_out(w320107));
	wire w360107;
	torch #(1'b1) c360107 (.i_clk(tick), .i_in(), .o_out(w360107));
	wire w400107;
	torch #(1'b1) c400107 (.i_clk(tick), .i_in(), .o_out(w400107));
	wire w440107;
	torch #(1'b1) c440107 (.i_clk(tick), .i_in(), .o_out(w440107));
	wire w530108;
	repeater #(1, 1'b0, 0, 0) c530108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530108));
	wire w1940110;

	wire w1950110;
	repeater #(1, 1'b0, 0, 0) c1950110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950110));
	wire w1960111;
	repeater #(1, 1'b0, 0, 0) c1960111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1960111));
	wire w1990111;
	repeater #(2, 1'b0, 0, 0) c1990111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990111));
	wire w1910112;
	repeater #(1, 1'b0, 0, 0) c1910112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910112));
	wire w2040112;
	repeater #(2, 1'b0, 0, 0) c2040112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040112));
	wire w1900113;
	assign outputs[57] = ();
	wire w1930113;

	wire w2020113;

	wire w1930114;

	wire w2020114;

	wire w1910115;
	repeater #(1, 1'b0, 0, 0) c1910115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910115));
	wire w2040115;
	repeater #(1, 1'b0, 0, 0) c2040115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040115));
	wire w250116;
	torch #(1'b1) c250116 (.i_clk(tick), .i_in(), .o_out(w250116));
	wire w290116;
	torch #(1'b1) c290116 (.i_clk(tick), .i_in(), .o_out(w290116));
	wire w330116;
	torch #(1'b1) c330116 (.i_clk(tick), .i_in(), .o_out(w330116));
	wire w370116;
	torch #(1'b1) c370116 (.i_clk(tick), .i_in(), .o_out(w370116));
	wire w410116;
	torch #(1'b1) c410116 (.i_clk(tick), .i_in(), .o_out(w410116));
	wire w450116;
	torch #(1'b1) c450116 (.i_clk(tick), .i_in(), .o_out(w450116));
	wire w490116;
	torch #(1'b1) c490116 (.i_clk(tick), .i_in(), .o_out(w490116));
	wire w260117;
	repeater #(1, 1'b0, 0, 0) c260117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260117));
	wire w300117;
	repeater #(1, 1'b0, 0, 0) c300117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300117));
	wire w340117;
	repeater #(1, 1'b0, 0, 0) c340117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340117));
	wire w380117;
	repeater #(1, 1'b1, 0, 0) c380117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380117));
	wire w420117;
	repeater #(1, 1'b0, 0, 0) c420117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420117));
	wire w460117;
	repeater #(1, 1'b0, 0, 0) c460117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460117));
	wire w500117;
	repeater #(1, 1'b0, 0, 0) c500117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500117));
	wire w240119;

	wire w260119;
	repeater #(1, 1'b0, 0, 0) c260119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260119));
	wire w280119;

	wire w300119;
	repeater #(1, 1'b0, 0, 0) c300119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300119));
	wire w320119;

	wire w340119;
	repeater #(1, 1'b0, 0, 0) c340119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340119));
	wire w360119;

	wire w380119;
	repeater #(1, 1'b1, 0, 0) c380119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380119));
	wire w400119;

	wire w420119;
	repeater #(1, 1'b0, 0, 0) c420119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420119));
	wire w440119;

	wire w460119;
	repeater #(1, 1'b0, 0, 0) c460119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460119));
	wire w480119;

	wire w500119;
	repeater #(1, 1'b0, 0, 0) c500119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500119));
	wire w320123;
	torch #(1'b1) c320123 (.i_clk(tick), .i_in(), .o_out(w320123));
	wire w360123;
	torch #(1'b1) c360123 (.i_clk(tick), .i_in(), .o_out(w360123));
	wire w400123;
	torch #(1'b1) c400123 (.i_clk(tick), .i_in(), .o_out(w400123));
	wire w440123;
	torch #(1'b1) c440123 (.i_clk(tick), .i_in(), .o_out(w440123));
	wire w530124;
	repeater #(1, 1'b0, 0, 0) c530124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530124));
	wire w250132;
	torch #(1'b1) c250132 (.i_clk(tick), .i_in(), .o_out(w250132));
	wire w290132;
	torch #(1'b1) c290132 (.i_clk(tick), .i_in(), .o_out(w290132));
	wire w330132;
	torch #(1'b1) c330132 (.i_clk(tick), .i_in(), .o_out(w330132));
	wire w370132;
	torch #(1'b0) c370132 (.i_clk(tick), .i_in(), .o_out(w370132));
	wire w410132;
	torch #(1'b1) c410132 (.i_clk(tick), .i_in(), .o_out(w410132));
	wire w450132;
	torch #(1'b1) c450132 (.i_clk(tick), .i_in(), .o_out(w450132));
	wire w490132;
	torch #(1'b1) c490132 (.i_clk(tick), .i_in(), .o_out(w490132));
	wire w260133;
	repeater #(1, 1'b0, 0, 0) c260133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260133));
	wire w300133;
	repeater #(1, 1'b0, 0, 0) c300133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300133));
	wire w340133;
	repeater #(1, 1'b0, 0, 0) c340133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340133));
	wire w380133;
	repeater #(1, 1'b1, 0, 0) c380133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380133));
	wire w420133;
	repeater #(1, 1'b0, 0, 0) c420133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420133));
	wire w460133;
	repeater #(1, 1'b0, 0, 0) c460133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460133));
	wire w500133;
	repeater #(1, 1'b0, 0, 0) c500133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500133));
	wire w240135;

	wire w260135;
	repeater #(1, 1'b0, 0, 0) c260135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260135));
	wire w280135;

	wire w300135;
	repeater #(1, 1'b0, 0, 0) c300135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300135));
	wire w320135;

	wire w340135;
	repeater #(1, 1'b0, 0, 0) c340135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340135));
	wire w360135;

	wire w380135;
	repeater #(1, 1'b1, 0, 0) c380135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380135));
	wire w400135;

	wire w420135;
	repeater #(1, 1'b0, 0, 0) c420135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420135));
	wire w440135;

	wire w460135;
	repeater #(1, 1'b0, 0, 0) c460135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460135));
	wire w480135;

	wire w500135;
	repeater #(1, 1'b0, 0, 0) c500135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500135));
	wire w250141;
	torch #(1'b1) c250141 (.i_clk(tick), .i_in(), .o_out(w250141));
	wire w290141;
	torch #(1'b1) c290141 (.i_clk(tick), .i_in(), .o_out(w290141));
	wire w330141;
	torch #(1'b1) c330141 (.i_clk(tick), .i_in(), .o_out(w330141));
	wire w370141;
	torch #(1'b0) c370141 (.i_clk(tick), .i_in(), .o_out(w370141));
	wire w410141;
	torch #(1'b1) c410141 (.i_clk(tick), .i_in(), .o_out(w410141));
	wire w450141;
	torch #(1'b1) c450141 (.i_clk(tick), .i_in(), .o_out(w450141));
	wire w490141;
	torch #(1'b1) c490141 (.i_clk(tick), .i_in(), .o_out(w490141));
	wire w260153;
	repeater #(1, 1'b0, 0, 0) c260153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260153));
	wire w300153;
	repeater #(1, 1'b0, 0, 0) c300153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300153));
	wire w340153;
	repeater #(1, 1'b0, 0, 0) c340153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340153));
	wire w380153;
	repeater #(1, 1'b1, 0, 0) c380153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380153));
	wire w420153;
	repeater #(1, 1'b0, 0, 0) c420153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420153));
	wire w460153;
	repeater #(1, 1'b0, 0, 0) c460153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460153));
	wire w500153;
	repeater #(1, 1'b0, 0, 0) c500153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500153));
	wire w250154;
	repeater #(1, 1'b1, 0, 0) c250154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250154));
	wire w290154;
	repeater #(1, 1'b1, 0, 0) c290154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290154));
	wire w330154;
	repeater #(1, 1'b1, 0, 0) c330154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330154));
	wire w370154;
	repeater #(1, 1'b1, 0, 0) c370154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w370154));
	wire w410154;
	repeater #(1, 1'b1, 0, 0) c410154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w410154));
	wire w450154;
	repeater #(1, 1'b1, 0, 0) c450154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w450154));
	wire w490154;
	repeater #(1, 1'b1, 0, 0) c490154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w490154));
	wire w280175;
	repeater #(1, 1'b0, 0, 0) c280175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w280175));
	wire w320175;
	repeater #(1, 1'b0, 0, 0) c320175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320175));
	wire w360175;
	repeater #(1, 1'b0, 0, 0) c360175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w360175));
	wire w400175;
	repeater #(1, 1'b0, 0, 0) c400175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400175));
	wire w440175;
	repeater #(1, 1'b0, 0, 0) c440175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w440175));
	wire w480175;
	repeater #(1, 1'b0, 0, 0) c480175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480175));
	wire w520175;
	repeater #(1, 1'b0, 0, 0) c520175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w520175));
	wire w2519;
	torch #(1'b1) c2519 (.i_clk(tick), .i_in(), .o_out(w2519));
	wire w2919;
	torch #(1'b1) c2919 (.i_clk(tick), .i_in(), .o_out(w2919));
	wire w3319;
	torch #(1'b1) c3319 (.i_clk(tick), .i_in(), .o_out(w3319));
	wire w3719;
	torch #(1'b0) c3719 (.i_clk(tick), .i_in(), .o_out(w3719));
	wire w4119;
	torch #(1'b1) c4119 (.i_clk(tick), .i_in(), .o_out(w4119));
	wire w4519;
	torch #(1'b1) c4519 (.i_clk(tick), .i_in(), .o_out(w4519));
	wire w4919;
	torch #(1'b1) c4919 (.i_clk(tick), .i_in(), .o_out(w4919));
	wire w141113;

	wire w175113;

	wire w1114;

	wire w35114;

	wire w140114;
	repeater #(1, 1'b1, 0, 0) c140114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140114));
	wire w174114;
	repeater #(1, 1'b1, 0, 0) c174114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174114));
	wire w0115;
	repeater #(1, 1'b1, 0, 0) c0115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0115));
	wire w34115;
	repeater #(1, 1'b1, 0, 0) c34115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34115));
	wire w139115;

	wire w173115;

	wire w207115;

	wire w33116;

	wire w138116;
	repeater #(1, 1'b1, 0, 0) c138116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138116));
	wire w172116;
	repeater #(1, 1'b1, 0, 0) c172116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172116));
	wire w206116;
	repeater #(1, 1'b1, 0, 0) c206116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206116));
	wire w32117;
	repeater #(1, 1'b1, 0, 0) c32117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32117));
	wire w137117;

	wire w171117;

	wire w205117;

	wire w31118;

	wire w136118;
	repeater #(1, 1'b1, 0, 0) c136118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136118));
	wire w170118;
	repeater #(1, 1'b1, 0, 0) c170118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170118));
	wire w204118;
	repeater #(1, 1'b1, 0, 0) c204118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204118));
	wire w30119;
	repeater #(1, 1'b1, 0, 0) c30119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30119));
	wire w135119;

	wire w169119;

	wire w203119;

	wire w29120;

	wire w134120;
	repeater #(1, 1'b1, 0, 0) c134120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134120));
	wire w168120;
	repeater #(1, 1'b1, 0, 0) c168120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168120));
	wire w202120;
	repeater #(1, 1'b1, 0, 0) c202120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202120));
	wire w28121;
	repeater #(1, 1'b1, 0, 0) c28121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28121));
	wire w133121;

	wire w167121;

	wire w201121;

	wire w27122;

	wire w132122;
	repeater #(1, 1'b1, 0, 0) c132122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132122));
	wire w166122;
	repeater #(1, 1'b1, 0, 0) c166122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166122));
	wire w200122;
	repeater #(1, 1'b1, 0, 0) c200122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200122));
	wire w26123;
	repeater #(1, 1'b1, 0, 0) c26123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26123));
	wire w131123;

	wire w165123;

	wire w199123;

	wire w25124;

	wire w130124;
	repeater #(1, 1'b1, 0, 0) c130124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130124));
	wire w164124;
	repeater #(1, 1'b1, 0, 0) c164124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164124));
	wire w198124;
	repeater #(1, 1'b1, 0, 0) c198124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198124));
	wire w24125;
	repeater #(1, 1'b1, 0, 0) c24125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24125));
	wire w129125;

	wire w163125;

	wire w197125;

	wire w23126;

	wire w128126;
	repeater #(1, 1'b1, 0, 0) c128126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128126));
	wire w162126;
	repeater #(1, 1'b1, 0, 0) c162126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162126));
	wire w196126;
	repeater #(1, 1'b1, 0, 0) c196126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196126));
	wire w22127;
	repeater #(1, 1'b1, 0, 0) c22127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22127));
	wire w127127;

	wire w161127;

	wire w195127;

	wire w21128;

	wire w126128;
	repeater #(1, 1'b0, 0, 0) c126128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126128));
	wire w160128;
	repeater #(1, 1'b0, 0, 0) c160128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160128));
	wire w194128;
	repeater #(1, 1'b0, 0, 0) c194128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194128));
	wire w20129;
	repeater #(1, 1'b0, 0, 0) c20129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20129));
	wire w125129;

	wire w159129;

	wire w193129;

	wire w19130;

	wire w124130;
	repeater #(1, 1'b1, 0, 0) c124130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124130));
	wire w158130;
	repeater #(1, 1'b1, 0, 0) c158130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158130));
	wire w192130;
	repeater #(1, 1'b1, 0, 0) c192130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192130));
	wire w18131;
	repeater #(1, 1'b1, 0, 0) c18131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18131));
	wire w123131;

	wire w157131;

	wire w191131;

	wire w17132;

	wire w122132;
	repeater #(1, 1'b1, 0, 0) c122132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122132));
	wire w156132;
	repeater #(1, 1'b1, 0, 0) c156132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156132));
	wire w190132;
	repeater #(1, 1'b1, 0, 0) c190132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190132));
	wire w16133;
	repeater #(1, 1'b1, 0, 0) c16133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16133));
	wire w121133;

	wire w155133;

	wire w189133;

	wire w15134;

	wire w120134;
	repeater #(1, 1'b1, 0, 0) c120134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120134));
	wire w154134;
	repeater #(1, 1'b1, 0, 0) c154134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154134));
	wire w188134;
	repeater #(1, 1'b1, 0, 0) c188134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188134));
	wire w14135;
	repeater #(1, 1'b1, 0, 0) c14135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14135));
	wire w119135;

	wire w153135;

	wire w187135;

	wire w13136;

	wire w56136;
	repeater #(1, 1'b1, 0, 0) c56136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56136));
	wire w118136;
	repeater #(1, 1'b1, 0, 0) c118136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118136));
	wire w152136;
	repeater #(1, 1'b1, 0, 0) c152136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152136));
	wire w186136;
	repeater #(1, 1'b1, 0, 0) c186136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186136));
	wire w12137;
	repeater #(1, 1'b1, 0, 0) c12137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12137));
	wire w117137;

	wire w151137;

	wire w185137;

	wire w11138;

	wire w116138;
	repeater #(1, 1'b1, 0, 0) c116138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116138));
	wire w150138;
	repeater #(1, 1'b1, 0, 0) c150138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150138));
	wire w184138;
	repeater #(1, 1'b1, 0, 0) c184138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184138));
	wire w10139;
	repeater #(1, 1'b1, 0, 0) c10139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10139));
	wire w115139;

	wire w149139;

	wire w183139;

	wire w9140;

	wire w114140;
	repeater #(1, 1'b1, 0, 0) c114140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114140));
	wire w148140;
	repeater #(1, 1'b1, 0, 0) c148140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148140));
	wire w182140;
	repeater #(1, 1'b1, 0, 0) c182140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182140));
	wire w8141;
	repeater #(1, 1'b1, 0, 0) c8141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8141));
	wire w165144;
	torch #(1'b0) c165144 (.i_clk(tick), .i_in(), .o_out(w165144));
	wire w169144;
	torch #(1'b0) c169144 (.i_clk(tick), .i_in(), .o_out(w169144));
	wire w173144;
	torch #(1'b0) c173144 (.i_clk(tick), .i_in(), .o_out(w173144));
	wire w177144;
	torch #(1'b1) c177144 (.i_clk(tick), .i_in(), .o_out(w177144));
	wire w181144;
	torch #(1'b0) c181144 (.i_clk(tick), .i_in(), .o_out(w181144));
	wire w185144;
	torch #(1'b0) c185144 (.i_clk(tick), .i_in(), .o_out(w185144));
	wire w189144;
	torch #(1'b0) c189144 (.i_clk(tick), .i_in(), .o_out(w189144));
	wire w201144;
	torch #(1'b0) c201144 (.i_clk(tick), .i_in(), .o_out(w201144));
	wire w205144;
	torch #(1'b0) c205144 (.i_clk(tick), .i_in(), .o_out(w205144));
	wire w1145;
	torch #(1'b1) c1145 (.i_clk(tick), .i_in(), .o_out(w1145));
	wire w5145;
	torch #(1'b1) c5145 (.i_clk(tick), .i_in(), .o_out(w5145));
	wire w9145;
	torch #(1'b1) c9145 (.i_clk(tick), .i_in(), .o_out(w9145));
	wire w13145;
	torch #(1'b0) c13145 (.i_clk(tick), .i_in(), .o_out(w13145));
	wire w17145;
	torch #(1'b0) c17145 (.i_clk(tick), .i_in(), .o_out(w17145));
	wire w112145;
	repeater #(2, 1'b1, 0, 0) c112145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112145));
	wire w146145;
	repeater #(2, 1'b1, 0, 0) c146145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146145));
	wire w24147;
	repeater #(1, 1'b1, 0, 0) c24147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24147));
	wire w28147;
	repeater #(1, 1'b1, 0, 0) c28147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28147));
	wire w32147;
	repeater #(1, 1'b1, 0, 0) c32147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32147));
	wire w36147;
	repeater #(1, 1'b0, 0, 0) c36147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36147));
	wire w40147;
	repeater #(1, 1'b1, 0, 0) c40147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40147));
	wire w44147;
	repeater #(1, 1'b1, 0, 0) c44147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44147));
	wire w48147;
	repeater #(1, 1'b1, 0, 0) c48147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48147));
	wire w98147;
	repeater #(1, 1'b1, 0, 0) c98147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98147));
	wire w104147;
	torch #(1'b1) c104147 (.i_clk(tick), .i_in(), .o_out(w104147));
	wire w114147;
	repeater #(1, 1'b1, 0, 0) c114147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114147));
	wire w120147;
	torch #(1'b1) c120147 (.i_clk(tick), .i_in(), .o_out(w120147));
	wire w132147;
	repeater #(1, 1'b1, 0, 0) c132147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132147));
	wire w138147;
	torch #(1'b1) c138147 (.i_clk(tick), .i_in(), .o_out(w138147));
	wire w148147;
	repeater #(1, 1'b1, 0, 0) c148147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148147));
	wire w154147;
	torch #(1'b1) c154147 (.i_clk(tick), .i_in(), .o_out(w154147));
	wire w24148;
	repeater #(1, 1'b1, 0, 0) c24148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24148));
	wire w26148;
	repeater #(1, 1'b0, 0, 0) c26148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26148));
	wire w28148;
	repeater #(1, 1'b1, 0, 0) c28148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28148));
	wire w30148;
	repeater #(1, 1'b0, 0, 0) c30148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30148));
	wire w32148;
	repeater #(1, 1'b1, 0, 0) c32148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32148));
	wire w34148;
	repeater #(1, 1'b0, 0, 0) c34148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34148));
	wire w36148;
	repeater #(1, 1'b0, 0, 0) c36148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36148));
	wire w38148;
	repeater #(1, 1'b0, 0, 0) c38148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38148));
	wire w40148;
	repeater #(1, 1'b1, 0, 0) c40148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40148));
	wire w42148;
	repeater #(1, 1'b0, 0, 0) c42148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42148));
	wire w44148;
	repeater #(1, 1'b1, 0, 0) c44148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44148));
	wire w46148;
	repeater #(1, 1'b0, 0, 0) c46148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46148));
	wire w48148;
	repeater #(1, 1'b1, 0, 0) c48148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48148));
	wire w50148;
	repeater #(1, 1'b0, 0, 0) c50148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50148));
	wire w25149;
	torch #(1'b0) c25149 (.i_clk(tick), .i_in(), .o_out(w25149));
	wire w29149;
	torch #(1'b0) c29149 (.i_clk(tick), .i_in(), .o_out(w29149));
	wire w33149;
	torch #(1'b0) c33149 (.i_clk(tick), .i_in(), .o_out(w33149));
	wire w37149;
	torch #(1'b0) c37149 (.i_clk(tick), .i_in(), .o_out(w37149));
	wire w41149;
	torch #(1'b0) c41149 (.i_clk(tick), .i_in(), .o_out(w41149));
	wire w45149;
	torch #(1'b0) c45149 (.i_clk(tick), .i_in(), .o_out(w45149));
	wire w49149;
	torch #(1'b0) c49149 (.i_clk(tick), .i_in(), .o_out(w49149));
	wire w105150;
	repeater #(1, 1'b1, 0, 0) c105150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105150));
	wire w121150;
	repeater #(1, 1'b1, 0, 0) c121150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121150));
	wire w139150;
	repeater #(1, 1'b1, 0, 0) c139150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139150));
	wire w155150;
	repeater #(1, 1'b1, 0, 0) c155150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155150));
	wire w98151;
	repeater #(1, 1'b1, 0, 0) c98151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98151));
	wire w114151;
	repeater #(1, 1'b1, 0, 0) c114151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114151));
	wire w132151;
	repeater #(1, 1'b1, 0, 0) c132151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132151));
	wire w148151;
	repeater #(1, 1'b1, 0, 0) c148151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148151));
	wire w165151;
	repeater #(1, 1'b1, 0, 0) c165151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165151));
	wire w169151;
	repeater #(1, 1'b1, 0, 0) c169151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169151));
	wire w173151;
	repeater #(1, 1'b1, 0, 0) c173151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173151));
	wire w177151;
	repeater #(1, 1'b0, 0, 0) c177151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177151));
	wire w181151;
	repeater #(1, 1'b1, 0, 0) c181151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181151));
	wire w185151;
	repeater #(1, 1'b1, 0, 0) c185151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185151));
	wire w189151;
	repeater #(1, 1'b1, 0, 0) c189151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189151));
	wire w201151;
	repeater #(1, 1'b1, 0, 0) c201151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201151));
	wire w205151;
	repeater #(1, 1'b1, 0, 0) c205151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205151));
	wire w1152;
	repeater #(1, 1'b0, 0, 0) c1152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1152));
	wire w5152;
	repeater #(1, 1'b0, 0, 0) c5152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5152));
	wire w9152;
	repeater #(1, 1'b0, 0, 0) c9152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9152));
	wire w13152;
	repeater #(1, 1'b1, 0, 0) c13152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13152));
	wire w17152;
	repeater #(1, 1'b1, 0, 0) c17152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17152));
	wire w103152;

	wire w119152;

	wire w137152;

	wire w153152;

	wire w111153;

	wire w145153;

	wire w98154;

	wire w108154;

	wire w113154;

	wire w114154;

	wire w132154;

	wire w142154;

	wire w147154;

	wire w148154;

	wire w171154;
	torch #(1'b0) c171154 (.i_clk(tick), .i_in(), .o_out(w171154));
	wire w175154;
	torch #(1'b0) c175154 (.i_clk(tick), .i_in(), .o_out(w175154));
	wire w179154;
	torch #(1'b1) c179154 (.i_clk(tick), .i_in(), .o_out(w179154));
	wire w183154;
	torch #(1'b1) c183154 (.i_clk(tick), .i_in(), .o_out(w183154));
	wire w207154;
	torch #(1'b0) c207154 (.i_clk(tick), .i_in(), .o_out(w207154));
	wire w3155;
	torch #(1'b0) c3155 (.i_clk(tick), .i_in(), .o_out(w3155));
	wire w7155;
	torch #(1'b0) c7155 (.i_clk(tick), .i_in(), .o_out(w7155));
	wire w11155;
	torch #(1'b0) c11155 (.i_clk(tick), .i_in(), .o_out(w11155));
	wire w32156;
	torch #(1'b1) c32156 (.i_clk(tick), .i_in(), .o_out(w32156));
	wire w36156;
	torch #(1'b1) c36156 (.i_clk(tick), .i_in(), .o_out(w36156));
	wire w40156;
	torch #(1'b1) c40156 (.i_clk(tick), .i_in(), .o_out(w40156));
	wire w44156;
	torch #(1'b1) c44156 (.i_clk(tick), .i_in(), .o_out(w44156));
	wire w106156;

	wire w140156;

	wire w97157;

	wire w112157;

	wire w113157;

	wire w131157;

	wire w146157;

	wire w147157;

	wire w98158;

	wire w102158;

	wire w106158;

	wire w132158;

	wire w136158;

	wire w140158;

	wire w26159;

	wire w30159;

	wire w34159;

	wire w38159;

	wire w42159;

	wire w46159;

	wire w50159;

	wire w122161;

	wire w156161;

	wire w95162;

	wire w96162;

	wire w99162;

	wire w100162;

	wire w103162;

	wire w104162;

	wire w107162;

	wire w108162;

	wire w111162;

	wire w112162;

	wire w115162;

	wire w116162;

	wire w119162;

	wire w120162;

	wire w129162;

	wire w130162;

	wire w133162;

	wire w134162;

	wire w137162;

	wire w138162;

	wire w141162;

	wire w142162;

	wire w145162;

	wire w146162;

	wire w149162;

	wire w150162;

	wire w153162;

	wire w154162;

	wire w93163;

	wire w127163;

	wire w108166;
	repeater #(1, 1'b1, 0, 0) c108166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108166));
	wire w112166;
	repeater #(1, 1'b1, 0, 0) c112166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112166));
	wire w116166;
	repeater #(1, 1'b0, 0, 0) c116166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116166));
	wire w142166;
	repeater #(1, 1'b1, 0, 0) c142166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142166));
	wire w146166;
	repeater #(1, 1'b1, 0, 0) c146166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146166));
	wire w150166;
	repeater #(1, 1'b1, 0, 0) c150166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150166));
	wire w94169;

	wire w98169;

	wire w114169;

	wire w118169;

	wire w128169;

	wire w132169;

	wire w148169;

	wire w152169;

	wire w166169;

	wire w167169;
	repeater #(1, 1'b1, 0, 0) c167169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167169));
	wire w171169;

	wire w172169;
	repeater #(1, 1'b1, 0, 0) c172169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172169));
	wire w176169;

	wire w177169;
	repeater #(1, 1'b1, 0, 0) c177169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177169));
	wire w5170;
	repeater #(1, 1'b1, 0, 0) c5170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5170));
	wire w6170;

	wire w10170;
	repeater #(1, 1'b1, 0, 0) c10170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10170));
	wire w11170;

	wire w15170;
	repeater #(1, 1'b1, 0, 0) c15170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15170));
	wire w16170;

	wire w26170;
	torch #(1'b0) c26170 (.i_clk(tick), .i_in(), .o_out(w26170));
	wire w30170;
	torch #(1'b0) c30170 (.i_clk(tick), .i_in(), .o_out(w30170));
	wire w34170;
	torch #(1'b0) c34170 (.i_clk(tick), .i_in(), .o_out(w34170));
	wire w38170;
	torch #(1'b1) c38170 (.i_clk(tick), .i_in(), .o_out(w38170));
	wire w42170;
	torch #(1'b0) c42170 (.i_clk(tick), .i_in(), .o_out(w42170));
	wire w46170;
	torch #(1'b0) c46170 (.i_clk(tick), .i_in(), .o_out(w46170));
	wire w50170;
	torch #(1'b0) c50170 (.i_clk(tick), .i_in(), .o_out(w50170));
	wire w96170;
	repeater #(1, 1'b1, 0, 0) c96170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96170));
	wire w130170;
	repeater #(1, 1'b1, 0, 0) c130170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130170));
	wire w90171;

	wire w103171;
	repeater #(1, 1'b1, 0, 0) c103171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103171));
	wire w124171;

	wire w137171;
	repeater #(1, 1'b1, 0, 0) c137171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137171));
	wire w32172;
	torch #(1'b1) c32172 (.i_clk(tick), .i_in(), .o_out(w32172));
	wire w36172;
	torch #(1'b1) c36172 (.i_clk(tick), .i_in(), .o_out(w36172));
	wire w40172;
	torch #(1'b1) c40172 (.i_clk(tick), .i_in(), .o_out(w40172));
	wire w44172;
	torch #(1'b1) c44172 (.i_clk(tick), .i_in(), .o_out(w44172));
	wire w58172;
	repeater #(1, 1'b1, 0, 0) c58172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58172));
	wire w60172;
	repeater #(1, 1'b1, 0, 0) c60172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60172));
	wire w62172;
	repeater #(1, 1'b1, 0, 0) c62172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62172));
	wire w98172;

	wire w114172;

	wire w132172;

	wire w148172;

	wire w90173;

	wire w106173;

	wire w124173;

	wire w140173;

	wire w166173;

	wire w167173;
	repeater #(1, 1'b0, 0, 0) c167173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167173));
	wire w171173;

	wire w172173;
	repeater #(1, 1'b0, 0, 0) c172173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172173));
	wire w176173;

	wire w177173;
	repeater #(1, 1'b1, 0, 0) c177173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177173));
	wire w5174;
	repeater #(1, 1'b1, 0, 0) c5174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5174));
	wire w6174;

	wire w10174;
	repeater #(1, 1'b0, 0, 0) c10174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10174));
	wire w11174;

	wire w15174;
	repeater #(1, 1'b1, 0, 0) c15174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15174));
	wire w16174;

	wire w93174;

	wire w101174;

	wire w103174;

	wire w104174;

	wire w109174;

	wire w117174;

	wire w127174;

	wire w135174;

	wire w137174;

	wire w138174;

	wire w143174;

	wire w151174;

	wire w26175;

	wire w30175;

	wire w34175;

	wire w38175;

	wire w42175;

	wire w46175;

	wire w50175;

	wire w95176;

	wire w96176;

	wire w111176;

	wire w112176;

	wire w129176;

	wire w130176;

	wire w145176;

	wire w146176;

	wire w186176;
	repeater #(1, 1'b1, 0, 0) c186176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186176));
	wire w204176;
	repeater #(1, 1'b1, 0, 0) c204176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204176));
	wire w166177;

	wire w167177;
	repeater #(1, 1'b0, 0, 0) c167177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167177));
	wire w171177;

	wire w172177;
	repeater #(1, 1'b0, 0, 0) c172177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172177));
	wire w176177;

	wire w177177;
	repeater #(1, 1'b0, 0, 0) c177177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177177));
	wire w5178;
	repeater #(1, 1'b1, 0, 0) c5178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5178));
	wire w6178;

	wire w10178;
	repeater #(1, 1'b0, 0, 0) c10178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10178));
	wire w11178;

	wire w15178;
	repeater #(1, 1'b0, 0, 0) c15178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15178));
	wire w16178;

	wire w101178;

	wire w103178;

	wire w104178;

	wire w117178;

	wire w135178;

	wire w137178;

	wire w138178;

	wire w151178;

	wire w194178;

	wire w193179;
	repeater #(1, 1'b1, 0, 0) c193179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193179));
	wire w98180;
	torch #(1'b1) c98180 (.i_clk(tick), .i_in(), .o_out(w98180));
	wire w99180;

	wire w114180;
	torch #(1'b1) c114180 (.i_clk(tick), .i_in(), .o_out(w114180));
	wire w115180;

	wire w132180;
	torch #(1'b1) c132180 (.i_clk(tick), .i_in(), .o_out(w132180));
	wire w133180;

	wire w148180;
	torch #(1'b1) c148180 (.i_clk(tick), .i_in(), .o_out(w148180));
	wire w149180;

	wire w99181;

	wire w101181;

	wire w115181;

	wire w117181;

	wire w133181;

	wire w135181;

	wire w149181;

	wire w151181;

	wire w165181;
	repeater #(1, 1'b1, 0, 0) c165181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165181));
	wire w197181;

	wire w17182;
	repeater #(1, 1'b0, 0, 0) c17182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17182));
	wire w169182;
	repeater #(1, 1'b0, 0, 0) c169182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169182));
	wire w194182;

	wire w13183;
	repeater #(1, 1'b0, 0, 0) c13183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13183));
	wire w101183;

	wire w102183;

	wire w103183;

	wire w117183;

	wire w118183;

	wire w119183;

	wire w135183;

	wire w136183;

	wire w137183;

	wire w151183;

	wire w152183;

	wire w153183;

	wire w175183;

	wire w179183;
	repeater #(1, 1'b0, 0, 0) c179183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179183));
	wire w193183;

	wire w195183;
	repeater #(2, 1'b1, 0, 0) c195183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195183));
	wire w198183;
	repeater #(2, 1'b0, 0, 0) c198183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198183));
	wire w3184;
	repeater #(1, 1'b1, 0, 0) c3184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3184));
	wire w7184;

	wire w96184;

	wire w97184;

	wire w103184;

	wire w112184;

	wire w113184;

	wire w119184;

	wire w130184;

	wire w131184;

	wire w137184;

	wire w146184;

	wire w147184;

	wire w153184;

	wire w176184;

	wire w182184;
	repeater #(2, 1'b1, 0, 0) c182184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182184));
	wire w185184;
	repeater #(2, 1'b0, 0, 0) c185184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185184));
	wire w187184;

	wire w203184;

	wire w205184;
	repeater #(2, 1'b0, 0, 0) c205184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205184));
	wire w0185;
	repeater #(2, 1'b1, 0, 0) c0185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0185));
	wire w6185;

	wire w175185;
	repeater #(2, 1'b0, 0, 0) c175185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175185));
	wire w186185;

	wire w204185;

	wire w7186;
	repeater #(2, 1'b1, 0, 0) c7186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7186));
	wire w26186;
	torch #(1'b0) c26186 (.i_clk(tick), .i_in(), .o_out(w26186));
	wire w30186;
	torch #(1'b0) c30186 (.i_clk(tick), .i_in(), .o_out(w30186));
	wire w34186;
	torch #(1'b0) c34186 (.i_clk(tick), .i_in(), .o_out(w34186));
	wire w38186;
	torch #(1'b1) c38186 (.i_clk(tick), .i_in(), .o_out(w38186));
	wire w42186;
	torch #(1'b0) c42186 (.i_clk(tick), .i_in(), .o_out(w42186));
	wire w46186;
	torch #(1'b0) c46186 (.i_clk(tick), .i_in(), .o_out(w46186));
	wire w50186;
	torch #(1'b0) c50186 (.i_clk(tick), .i_in(), .o_out(w50186));
	wire w101186;
	repeater #(1, 1'b0, 0, 0) c101186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101186));
	wire w103186;
	torch #(1'b0) c103186 (.i_clk(tick), .i_in(), .o_out(w103186));
	wire w109186;
	torch #(1'b0) c109186 (.i_clk(tick), .i_in(), .o_out(w109186));
	wire w117186;
	repeater #(1, 1'b0, 0, 0) c117186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117186));
	wire w119186;
	torch #(1'b0) c119186 (.i_clk(tick), .i_in(), .o_out(w119186));
	wire w135186;
	repeater #(1, 1'b0, 0, 0) c135186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135186));
	wire w137186;
	torch #(1'b0) c137186 (.i_clk(tick), .i_in(), .o_out(w137186));
	wire w143186;
	torch #(1'b0) c143186 (.i_clk(tick), .i_in(), .o_out(w143186));
	wire w151186;
	repeater #(1, 1'b0, 0, 0) c151186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151186));
	wire w153186;
	torch #(1'b0) c153186 (.i_clk(tick), .i_in(), .o_out(w153186));
	wire w169186;

	wire w170186;

	wire w183186;

	wire w207186;

	wire w12187;

	wire w13187;

	wire w168187;

	wire w177187;

	wire w5188;

	wire w14188;

	wire w32188;
	torch #(1'b1) c32188 (.i_clk(tick), .i_in(), .o_out(w32188));
	wire w36188;
	torch #(1'b1) c36188 (.i_clk(tick), .i_in(), .o_out(w36188));
	wire w40188;
	torch #(1'b1) c40188 (.i_clk(tick), .i_in(), .o_out(w40188));
	wire w44188;
	torch #(1'b1) c44188 (.i_clk(tick), .i_in(), .o_out(w44188));
	wire w105188;
	repeater #(1, 1'b1, 0, 0) c105188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105188));
	wire w121188;
	repeater #(1, 1'b1, 0, 0) c121188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121188));
	wire w139188;
	repeater #(1, 1'b1, 0, 0) c139188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139188));
	wire w155188;
	repeater #(1, 1'b1, 0, 0) c155188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155188));
	wire w171188;

	wire w201188;
	assign outputs[58] = ();
	wire w11189;

	wire w102190;
	torch #(1'b1) c102190 (.i_clk(tick), .i_in(), .o_out(w102190));
	wire w118190;
	torch #(1'b1) c118190 (.i_clk(tick), .i_in(), .o_out(w118190));
	wire w136190;
	torch #(1'b1) c136190 (.i_clk(tick), .i_in(), .o_out(w136190));
	wire w152190;
	torch #(1'b1) c152190 (.i_clk(tick), .i_in(), .o_out(w152190));
	wire w26191;

	wire w30191;

	wire w34191;

	wire w38191;

	wire w42191;

	wire w46191;

	wire w50191;

	wire w110192;
	torch #(1'b1) c110192 (.i_clk(tick), .i_in(), .o_out(w110192));
	wire w144192;
	torch #(1'b1) c144192 (.i_clk(tick), .i_in(), .o_out(w144192));
	wire w101193;
	repeater #(2, 1'b0, 0, 0) c101193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101193));
	wire w117193;
	repeater #(2, 1'b0, 0, 0) c117193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117193));
	wire w135193;
	repeater #(2, 1'b0, 0, 0) c135193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135193));
	wire w151193;
	repeater #(2, 1'b0, 0, 0) c151193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151193));
	wire w111194;
	repeater #(2, 1'b0, 0, 0) c111194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111194));
	wire w145194;
	repeater #(2, 1'b0, 0, 0) c145194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145194));
	wire w121196;
	repeater #(1, 1'b0, 0, 0) c121196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121196));
	wire w155196;
	repeater #(1, 1'b0, 0, 0) c155196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155196));
	wire w123197;
	repeater #(1, 1'b0, 0, 0) c123197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123197));
	wire w157197;
	repeater #(1, 1'b0, 0, 0) c157197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157197));
	wire w261102;
	torch #(1'b0) c261102 (.i_clk(tick), .i_in(), .o_out(w261102));
	wire w301102;
	torch #(1'b0) c301102 (.i_clk(tick), .i_in(), .o_out(w301102));
	wire w341102;
	torch #(1'b0) c341102 (.i_clk(tick), .i_in(), .o_out(w341102));
	wire w381102;
	torch #(1'b1) c381102 (.i_clk(tick), .i_in(), .o_out(w381102));
	wire w421102;
	torch #(1'b0) c421102 (.i_clk(tick), .i_in(), .o_out(w421102));
	wire w461102;
	torch #(1'b0) c461102 (.i_clk(tick), .i_in(), .o_out(w461102));
	wire w501102;
	torch #(1'b0) c501102 (.i_clk(tick), .i_in(), .o_out(w501102));
	wire w321104;
	torch #(1'b1) c321104 (.i_clk(tick), .i_in(), .o_out(w321104));
	wire w361104;
	torch #(1'b1) c361104 (.i_clk(tick), .i_in(), .o_out(w361104));
	wire w401104;
	torch #(1'b1) c401104 (.i_clk(tick), .i_in(), .o_out(w401104));
	wire w441104;
	torch #(1'b1) c441104 (.i_clk(tick), .i_in(), .o_out(w441104));
	wire w261107;

	wire w301107;

	wire w341107;

	wire w381107;

	wire w421107;

	wire w461107;

	wire w501107;

	wire w1881110;

	wire w2061110;

	wire w261118;
	torch #(1'b0) c261118 (.i_clk(tick), .i_in(), .o_out(w261118));
	wire w301118;
	torch #(1'b0) c301118 (.i_clk(tick), .i_in(), .o_out(w301118));
	wire w341118;
	torch #(1'b0) c341118 (.i_clk(tick), .i_in(), .o_out(w341118));
	wire w381118;
	torch #(1'b1) c381118 (.i_clk(tick), .i_in(), .o_out(w381118));
	wire w421118;
	torch #(1'b0) c421118 (.i_clk(tick), .i_in(), .o_out(w421118));
	wire w461118;
	torch #(1'b0) c461118 (.i_clk(tick), .i_in(), .o_out(w461118));
	wire w501118;
	torch #(1'b0) c501118 (.i_clk(tick), .i_in(), .o_out(w501118));
	wire w321120;
	torch #(1'b1) c321120 (.i_clk(tick), .i_in(), .o_out(w321120));
	wire w361120;
	torch #(1'b1) c361120 (.i_clk(tick), .i_in(), .o_out(w361120));
	wire w401120;
	torch #(1'b1) c401120 (.i_clk(tick), .i_in(), .o_out(w401120));
	wire w441120;
	torch #(1'b1) c441120 (.i_clk(tick), .i_in(), .o_out(w441120));
	wire w261123;

	wire w301123;

	wire w341123;

	wire w381123;

	wire w421123;

	wire w461123;

	wire w501123;

	wire w261134;
	torch #(1'b0) c261134 (.i_clk(tick), .i_in(), .o_out(w261134));
	wire w301134;
	torch #(1'b0) c301134 (.i_clk(tick), .i_in(), .o_out(w301134));
	wire w341134;
	torch #(1'b0) c341134 (.i_clk(tick), .i_in(), .o_out(w341134));
	wire w381134;
	torch #(1'b1) c381134 (.i_clk(tick), .i_in(), .o_out(w381134));
	wire w421134;
	torch #(1'b0) c421134 (.i_clk(tick), .i_in(), .o_out(w421134));
	wire w461134;
	torch #(1'b0) c461134 (.i_clk(tick), .i_in(), .o_out(w461134));
	wire w501134;
	torch #(1'b0) c501134 (.i_clk(tick), .i_in(), .o_out(w501134));
	wire w801;
	assign outputs[59] = ();
	wire w1001;
	assign outputs[60] = ();
	wire w1201;
	assign outputs[61] = ();
	wire w1401;
	assign outputs[62] = ();
	wire w1601;
	assign outputs[63] = ();
	wire w1801;
	assign outputs[64] = ();
	wire w2001;
	assign outputs[65] = ();
	wire w2201;
	assign outputs[66] = ();
	wire w2401;
	assign outputs[67] = ();
	wire w2601;
	assign outputs[68] = ();
	wire w2801;
	assign outputs[69] = ();
	wire w3001;
	assign outputs[70] = ();
	wire w3201;
	assign outputs[71] = ();
	wire w3401;
	assign outputs[72] = ();
	wire w802;
	repeater #(1, 1'b0, 0, 0) c802 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w802));
	wire w1002;
	repeater #(1, 1'b0, 0, 0) c1002 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1002));
	wire w1202;
	repeater #(1, 1'b0, 0, 0) c1202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1202));
	wire w1402;
	repeater #(1, 1'b0, 0, 0) c1402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1402));
	wire w1602;
	repeater #(1, 1'b0, 0, 0) c1602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1602));
	wire w1802;
	repeater #(1, 1'b0, 0, 0) c1802 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1802));
	wire w2002;
	repeater #(1, 1'b0, 0, 0) c2002 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2002));
	wire w2202;
	repeater #(1, 1'b1, 0, 0) c2202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2202));
	wire w2402;
	repeater #(1, 1'b0, 0, 0) c2402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2402));
	wire w2602;
	repeater #(1, 1'b0, 0, 0) c2602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2602));
	wire w2802;
	repeater #(1, 1'b0, 0, 0) c2802 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2802));
	wire w3002;
	repeater #(1, 1'b0, 0, 0) c3002 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3002));
	wire w3202;
	repeater #(1, 1'b0, 0, 0) c3202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3202));
	wire w3402;
	repeater #(1, 1'b0, 0, 0) c3402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3402));
	wire w909;
	repeater #(2, 1'b1, 0, 0) c909 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w909));
	wire w1309;
	repeater #(2, 1'b1, 0, 0) c1309 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1309));
	wire w1709;
	repeater #(2, 1'b1, 0, 0) c1709 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1709));
	wire w2109;
	repeater #(2, 1'b0, 0, 0) c2109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2109));
	wire w2509;
	repeater #(2, 1'b1, 0, 0) c2509 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2509));
	wire w2909;
	repeater #(2, 1'b1, 0, 0) c2909 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2909));
	wire w3309;
	repeater #(2, 1'b1, 0, 0) c3309 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3309));
	wire w7014;
	repeater #(1, 1'b1, 0, 0) c7014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7014));
	wire w11014;
	repeater #(1, 1'b1, 0, 0) c11014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11014));
	wire w15014;
	repeater #(1, 1'b1, 0, 0) c15014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15014));
	wire w19014;
	repeater #(1, 1'b0, 0, 0) c19014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19014));
	wire w23014;
	repeater #(1, 1'b1, 0, 0) c23014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23014));
	wire w27014;
	repeater #(1, 1'b1, 0, 0) c27014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27014));
	wire w31014;
	repeater #(1, 1'b1, 0, 0) c31014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31014));
	wire w9015;

	wire w13015;

	wire w17015;

	wire w21015;

	wire w25015;

	wire w29015;

	wire w33015;

	wire w8016;

	wire w12016;

	wire w16016;

	wire w20016;

	wire w24016;

	wire w28016;

	wire w32016;

	wire w9017;
	torch #(1'b1) c9017 (.i_clk(tick), .i_in(), .o_out(w9017));
	wire w13017;
	torch #(1'b1) c13017 (.i_clk(tick), .i_in(), .o_out(w13017));
	wire w17017;
	torch #(1'b1) c17017 (.i_clk(tick), .i_in(), .o_out(w17017));
	wire w21017;
	torch #(1'b1) c21017 (.i_clk(tick), .i_in(), .o_out(w21017));
	wire w25017;
	torch #(1'b1) c25017 (.i_clk(tick), .i_in(), .o_out(w25017));
	wire w29017;
	torch #(1'b1) c29017 (.i_clk(tick), .i_in(), .o_out(w29017));
	wire w33017;
	torch #(1'b1) c33017 (.i_clk(tick), .i_in(), .o_out(w33017));
	wire w7018;
	repeater #(1, 1'b1, 0, 0) c7018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7018));
	wire w11018;
	repeater #(1, 1'b1, 0, 0) c11018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11018));
	wire w15018;
	repeater #(1, 1'b1, 0, 0) c15018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15018));
	wire w19018;
	repeater #(1, 1'b1, 0, 0) c19018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19018));
	wire w23018;
	repeater #(1, 1'b1, 0, 0) c23018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23018));
	wire w27018;
	repeater #(1, 1'b1, 0, 0) c27018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w27018));
	wire w31018;
	repeater #(1, 1'b1, 0, 0) c31018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31018));
	wire w34076;

	wire w32078;

	wire w30080;

	wire w28082;

	wire w26084;

	wire w92088;
	repeater #(2, 1'b1, 0, 0) c92088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92088));
	wire w126088;
	repeater #(2, 1'b1, 0, 0) c126088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126088));
	wire w9090;
	torch #(1'b1) c9090 (.i_clk(tick), .i_in(), .o_out(w9090));
	wire w13090;
	torch #(1'b1) c13090 (.i_clk(tick), .i_in(), .o_out(w13090));
	wire w17090;
	torch #(1'b1) c17090 (.i_clk(tick), .i_in(), .o_out(w17090));
	wire w21090;
	torch #(1'b1) c21090 (.i_clk(tick), .i_in(), .o_out(w21090));
	wire w25090;
	torch #(1'b1) c25090 (.i_clk(tick), .i_in(), .o_out(w25090));
	wire w29090;
	torch #(1'b1) c29090 (.i_clk(tick), .i_in(), .o_out(w29090));
	wire w33090;
	torch #(1'b1) c33090 (.i_clk(tick), .i_in(), .o_out(w33090));
	wire w84090;
	torch #(1'b1) c84090 (.i_clk(tick), .i_in(), .o_out(w84090));
	wire w94090;
	repeater #(1, 1'b1, 0, 0) c94090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94090));
	wire w100090;
	torch #(1'b1) c100090 (.i_clk(tick), .i_in(), .o_out(w100090));
	wire w118090;
	torch #(1'b1) c118090 (.i_clk(tick), .i_in(), .o_out(w118090));
	wire w128090;
	repeater #(1, 1'b1, 0, 0) c128090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128090));
	wire w134090;
	torch #(1'b1) c134090 (.i_clk(tick), .i_in(), .o_out(w134090));
	wire w10093;
	repeater #(2, 1'b0, 0, 0) c10093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10093));
	wire w14093;
	repeater #(2, 1'b0, 0, 0) c14093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14093));
	wire w18093;
	repeater #(2, 1'b0, 0, 0) c18093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18093));
	wire w22093;
	repeater #(2, 1'b0, 0, 0) c22093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22093));
	wire w26093;
	repeater #(1, 1'b0, 0, 0) c26093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26093));
	wire w30093;
	repeater #(1, 1'b0, 0, 0) c30093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30093));
	wire w34093;
	repeater #(1, 1'b0, 0, 0) c34093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34093));
	wire w101093;
	repeater #(1, 1'b1, 0, 0) c101093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101093));
	wire w135093;
	repeater #(1, 1'b1, 0, 0) c135093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135093));
	wire w23094;
	repeater #(1, 1'b0, 0, 0) c23094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23094));
	wire w35094;
	repeater #(2, 1'b0, 0, 0) c35094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35094));
	wire w94094;
	repeater #(1, 1'b1, 0, 0) c94094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94094));
	wire w107094;

	wire w128094;
	repeater #(1, 1'b1, 0, 0) c128094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128094));
	wire w141094;

	wire w83095;

	wire w99095;

	wire w117095;

	wire w133095;

	wire w91096;

	wire w107096;

	wire w125096;

	wire w141096;

	wire w88097;

	wire w93097;

	wire w94097;

	wire w104097;

	wire w122097;

	wire w127097;

	wire w128097;

	wire w138097;

	wire w6099;
	repeater #(1, 1'b0, 0, 0) c6099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6099));
	wire w12099;
	repeater #(1, 1'b0, 0, 0) c12099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12099));
	wire w32099;
	repeater #(1, 1'b0, 0, 0) c32099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32099));
	wire w86099;

	wire w102099;

	wire w120099;

	wire w136099;

	wire w920100;

	wire w930100;

	wire w1260100;

	wire w1270100;

	wire w780101;

	wire w1120101;

	wire w1550101;
	repeater #(2, 1'b1, 0, 0) c1550101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550101));
	wire w1570101;
	repeater #(1, 1'b1, 0, 0) c1570101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570101));
	wire w1590101;
	repeater #(2, 1'b1, 0, 0) c1590101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1590101));
	wire w1610101;
	repeater #(1, 1'b0, 0, 0) c1610101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610101));
	wire w1630101;
	repeater #(2, 1'b0, 0, 0) c1630101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630101));
	wire w1650101;
	repeater #(1, 1'b1, 0, 0) c1650101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1650101));
	wire w1670101;
	repeater #(2, 1'b0, 0, 0) c1670101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1670101));
	wire w1690101;
	repeater #(1, 1'b1, 0, 0) c1690101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1690101));
	wire w1890101;
	repeater #(1, 1'b1, 0, 0) c1890101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1890101));
	wire w1910101;
	repeater #(2, 1'b1, 0, 0) c1910101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910101));
	wire w1930101;
	repeater #(1, 1'b0, 0, 0) c1930101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1930101));
	wire w1950101;
	repeater #(2, 1'b1, 0, 0) c1950101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950101));
	wire w1970101;
	repeater #(1, 1'b0, 0, 0) c1970101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970101));
	wire w1990101;
	repeater #(2, 1'b1, 0, 0) c1990101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990101));
	wire w2010101;
	repeater #(1, 1'b0, 0, 0) c2010101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010101));
	wire w2030101;
	repeater #(2, 1'b1, 0, 0) c2030101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030101));
	wire w790103;
	repeater #(1, 1'b1, 0, 0) c790103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w790103));
	wire w830103;
	repeater #(1, 1'b1, 0, 0) c830103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w830103));
	wire w870103;
	repeater #(1, 1'b1, 0, 0) c870103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w870103));
	wire w910103;
	repeater #(1, 1'b1, 0, 0) c910103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w910103));
	wire w950103;
	repeater #(1, 1'b1, 0, 0) c950103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w950103));
	wire w990103;
	repeater #(1, 1'b1, 0, 0) c990103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990103));
	wire w1030103;
	repeater #(1, 1'b0, 0, 0) c1030103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030103));
	wire w1130103;
	repeater #(1, 1'b1, 0, 0) c1130103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1130103));
	wire w1170103;
	repeater #(1, 1'b1, 0, 0) c1170103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1170103));
	wire w1210103;
	repeater #(1, 1'b1, 0, 0) c1210103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1210103));
	wire w1250103;
	repeater #(1, 1'b1, 0, 0) c1250103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1250103));
	wire w1290103;
	repeater #(1, 1'b1, 0, 0) c1290103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1290103));
	wire w1330103;
	repeater #(1, 1'b1, 0, 0) c1330103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1330103));
	wire w1370103;
	repeater #(1, 1'b1, 0, 0) c1370103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370103));
	wire w1640103;

	wire w1940103;

	wire w1560104;

	wire w1600104;

	wire w1630104;

	wire w1650104;

	wire w1680104;

	wire w1900104;

	wire w1930104;

	wire w1950104;

	wire w1980104;

	wire w2020104;

	wire w1550105;

	wire w1570105;

	wire w1590105;

	wire w1610105;

	wire w1640105;

	wire w1670105;

	wire w1690105;

	wire w1890105;

	wire w1910105;

	wire w1940105;

	wire w1970105;

	wire w1990105;

	wire w2010105;

	wire w2030105;

	wire w1600106;

	wire w1980106;

	wire w80107;
	torch #(1'b1) c80107 (.i_clk(tick), .i_in(), .o_out(w80107));
	wire w120107;
	torch #(1'b1) c120107 (.i_clk(tick), .i_in(), .o_out(w120107));
	wire w160107;
	torch #(1'b1) c160107 (.i_clk(tick), .i_in(), .o_out(w160107));
	wire w200107;
	torch #(1'b1) c200107 (.i_clk(tick), .i_in(), .o_out(w200107));
	wire w240107;
	torch #(1'b1) c240107 (.i_clk(tick), .i_in(), .o_out(w240107));
	wire w280107;
	torch #(1'b1) c280107 (.i_clk(tick), .i_in(), .o_out(w280107));
	wire w320107;
	torch #(1'b1) c320107 (.i_clk(tick), .i_in(), .o_out(w320107));
	wire w1560107;

	wire w1600107;

	wire w1610107;

	wire w1650107;

	wire w1670107;

	wire w1690107;

	wire w1890107;

	wire w1910107;

	wire w1930107;

	wire w1970107;

	wire w1980107;

	wire w2020107;

	wire w1620108;

	wire w1960108;

	wire w1530109;

	wire w1580109;

	wire w1590109;

	wire w1990109;

	wire w2000109;

	wire w2050109;

	wire w1510110;
	repeater #(1, 1'b1, 0, 0) c1510110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510110));
	wire w1560110;
	repeater #(1, 1'b1, 0, 0) c1560110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560110));
	wire w2020110;
	repeater #(1, 1'b1, 0, 0) c2020110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020110));
	wire w2070110;
	repeater #(1, 1'b1, 0, 0) c2070110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070110));
	wire w1610111;
	repeater #(1, 1'b1, 0, 0) c1610111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610111));
	wire w1970111;
	repeater #(1, 1'b1, 0, 0) c1970111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970111));
	wire w860112;

	wire w1200112;

	wire w840113;
	repeater #(1, 1'b1, 0, 0) c840113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840113));
	wire w1180113;
	repeater #(1, 1'b1, 0, 0) c1180113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1180113));
	wire w750114;
	repeater #(1, 1'b1, 0, 0) c750114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w750114));
	wire w780114;

	wire w910114;
	repeater #(1, 1'b1, 0, 0) c910114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w910114));
	wire w1090114;
	repeater #(1, 1'b1, 0, 0) c1090114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1090114));
	wire w1120114;

	wire w1250114;
	repeater #(1, 1'b1, 0, 0) c1250114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1250114));
	wire w1510114;
	repeater #(1, 1'b1, 0, 0) c1510114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510114));
	wire w1560114;
	repeater #(1, 1'b1, 0, 0) c1560114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560114));
	wire w1610114;
	repeater #(1, 1'b1, 0, 0) c1610114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610114));
	wire w1970114;
	repeater #(1, 1'b1, 0, 0) c1970114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970114));
	wire w2020114;
	repeater #(1, 1'b1, 0, 0) c2020114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020114));
	wire w2070114;
	repeater #(1, 1'b1, 0, 0) c2070114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070114));
	wire w60115;
	repeater #(1, 1'b0, 0, 0) c60115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60115));
	wire w120115;
	repeater #(1, 1'b0, 0, 0) c120115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120115));
	wire w320115;
	repeater #(1, 1'b0, 0, 0) c320115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320115));
	wire w860115;

	wire w1020115;

	wire w1200115;

	wire w1360115;

	wire w780116;

	wire w1120116;

	wire w750117;

	wire w760117;

	wire w810117;

	wire w890117;

	wire w910117;

	wire w920117;

	wire w1050117;

	wire w1090117;

	wire w1100117;

	wire w1150117;

	wire w1230117;

	wire w1250117;

	wire w1260117;

	wire w1390117;

	wire w1510118;
	repeater #(1, 1'b0, 0, 0) c1510118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510118));
	wire w1560118;
	repeater #(1, 1'b0, 0, 0) c1560118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560118));
	wire w1610118;
	repeater #(1, 1'b1, 0, 0) c1610118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610118));
	wire w1970118;
	repeater #(1, 1'b1, 0, 0) c1970118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970118));
	wire w2020118;
	repeater #(1, 1'b0, 0, 0) c2020118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020118));
	wire w2070118;
	repeater #(1, 1'b0, 0, 0) c2070118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070118));
	wire w830119;

	wire w840119;

	wire w990119;

	wire w1170119;

	wire w1180119;

	wire w1330119;

	wire w750121;

	wire w760121;

	wire w890121;

	wire w910121;

	wire w920121;

	wire w1050121;

	wire w1090121;

	wire w1100121;

	wire w1230121;

	wire w1250121;

	wire w1260121;

	wire w1390121;

	wire w1770121;

	wire w1510122;
	repeater #(2, 1'b0, 0, 0) c1510122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510122));
	wire w1560122;
	repeater #(2, 1'b0, 0, 0) c1560122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560122));
	wire w1610122;
	repeater #(2, 1'b0, 0, 0) c1610122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610122));
	wire w1970122;
	repeater #(2, 1'b0, 0, 0) c1970122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970122));
	wire w2020122;
	repeater #(2, 1'b0, 0, 0) c2020122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020122));
	wire w2070122;
	repeater #(2, 1'b0, 0, 0) c2070122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070122));
	wire w80123;
	torch #(1'b1) c80123 (.i_clk(tick), .i_in(), .o_out(w80123));
	wire w120123;
	torch #(1'b1) c120123 (.i_clk(tick), .i_in(), .o_out(w120123));
	wire w160123;
	torch #(1'b1) c160123 (.i_clk(tick), .i_in(), .o_out(w160123));
	wire w200123;
	torch #(1'b1) c200123 (.i_clk(tick), .i_in(), .o_out(w200123));
	wire w240123;
	torch #(1'b1) c240123 (.i_clk(tick), .i_in(), .o_out(w240123));
	wire w280123;
	torch #(1'b1) c280123 (.i_clk(tick), .i_in(), .o_out(w280123));
	wire w320123;
	torch #(1'b1) c320123 (.i_clk(tick), .i_in(), .o_out(w320123));
	wire w860123;
	torch #(1'b1) c860123 (.i_clk(tick), .i_in(), .o_out(w860123));
	wire w870123;

	wire w1020123;
	torch #(1'b1) c1020123 (.i_clk(tick), .i_in(), .o_out(w1020123));
	wire w1030123;

	wire w1200123;
	torch #(1'b1) c1200123 (.i_clk(tick), .i_in(), .o_out(w1200123));
	wire w1210123;

	wire w1360123;
	torch #(1'b1) c1360123 (.i_clk(tick), .i_in(), .o_out(w1360123));
	wire w1370123;

	wire w1520123;
	repeater #(2, 1'b1, 0, 0) c1520123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520123));
	wire w1790123;

	wire w2060123;
	repeater #(2, 1'b1, 0, 0) c2060123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060123));
	wire w870124;

	wire w890124;

	wire w1030124;

	wire w1050124;

	wire w1210124;

	wire w1230124;

	wire w1370124;

	wire w1390124;

	wire w1500124;

	wire w1510124;

	wire w1570124;
	repeater #(1, 1'b1, 0, 0) c1570124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570124));
	wire w1580124;
	repeater #(2, 1'b1, 0, 0) c1580124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580124));
	wire w1800124;

	wire w2000124;
	repeater #(2, 1'b0, 0, 0) c2000124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2000124));
	wire w2010124;
	repeater #(1, 1'b0, 0, 0) c2010124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010124));
	wire w2070124;

	wire w00125;

	wire w1540125;
	repeater #(2, 1'b1, 0, 0) c1540125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540125));
	wire w1550125;
	repeater #(2, 1'b1, 0, 0) c1550125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550125));
	wire w1570125;

	wire w1710125;
	repeater #(1, 1'b0, 0, 0) c1710125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710125));
	wire w1720125;

	wire w1800125;
	repeater #(1, 1'b1, 0, 0) c1800125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800125));
	wire w1860125;

	wire w1870125;
	repeater #(1, 1'b0, 0, 0) c1870125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870125));
	wire w2010125;

	wire w2030125;
	repeater #(2, 1'b0, 0, 0) c2030125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030125));
	wire w2040125;
	repeater #(2, 1'b0, 0, 0) c2040125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040125));
	wire w890126;

	wire w900126;

	wire w910126;

	wire w1050126;

	wire w1060126;

	wire w1070126;

	wire w1230126;

	wire w1240126;

	wire w1250126;

	wire w1390126;

	wire w1400126;

	wire w1410126;

	wire w1550126;

	wire w1570126;
	repeater #(1, 1'b1, 0, 0) c1570126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570126));
	wire w1680126;

	wire w1690126;

	wire w1890126;

	wire w1900126;

	wire w2010126;
	repeater #(1, 1'b1, 0, 0) c2010126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010126));
	wire w2030126;

	wire w840127;

	wire w850127;

	wire w910127;

	wire w1000127;

	wire w1010127;

	wire w1070127;

	wire w1180127;

	wire w1190127;

	wire w1250127;

	wire w1340127;

	wire w1350127;

	wire w1410127;

	wire w1510127;

	wire w1550127;

	wire w1790127;

	wire w1800127;

	wire w2030127;

	wire w2070127;

	wire w1510128;

	wire w1530128;
	repeater #(1, 1'b0, 0, 0) c1530128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1530128));
	wire w1580128;

	wire w1620128;

	wire w1680128;
	repeater #(1, 1'b0, 0, 0) c1680128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1680128));
	wire w1760128;

	wire w1770128;
	repeater #(1, 1'b1, 0, 0) c1770128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770128));
	wire w1900128;
	repeater #(1, 1'b0, 0, 0) c1900128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1900128));
	wire w1960128;

	wire w2000128;

	wire w2050128;
	repeater #(1, 1'b1, 0, 0) c2050128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2050128));
	wire w2070128;

	wire w890129;
	repeater #(1, 1'b0, 0, 0) c890129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w890129));
	wire w910129;
	torch #(1'b0) c910129 (.i_clk(tick), .i_in(), .o_out(w910129));
	wire w970129;
	torch #(1'b0) c970129 (.i_clk(tick), .i_in(), .o_out(w970129));
	wire w1050129;
	repeater #(1, 1'b1, 0, 0) c1050129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1050129));
	wire w1070129;
	torch #(1'b0) c1070129 (.i_clk(tick), .i_in(), .o_out(w1070129));
	wire w1230129;
	repeater #(1, 1'b0, 0, 0) c1230129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230129));
	wire w1250129;
	torch #(1'b0) c1250129 (.i_clk(tick), .i_in(), .o_out(w1250129));
	wire w1310129;
	torch #(1'b0) c1310129 (.i_clk(tick), .i_in(), .o_out(w1310129));
	wire w1390129;
	repeater #(1, 1'b1, 0, 0) c1390129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390129));
	wire w1410129;
	torch #(1'b0) c1410129 (.i_clk(tick), .i_in(), .o_out(w1410129));
	wire w1580129;

	wire w1600129;
	repeater #(1, 1'b0, 0, 0) c1600129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1600129));
	wire w1610129;

	wire w1680129;

	wire w1850129;

	wire w1900129;

	wire w1970129;

	wire w1980129;
	repeater #(1, 1'b1, 0, 0) c1980129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980129));
	wire w2000129;

	wire w1540130;

	wire w1690130;

	wire w1730130;
	repeater #(1, 1'b1, 0, 0) c1730130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1730130));
	wire w1860130;
	repeater #(2, 1'b1, 0, 0) c1860130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860130));
	wire w1890130;

	wire w2040130;

	wire w60131;
	repeater #(1, 1'b0, 0, 0) c60131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60131));
	wire w120131;
	repeater #(1, 1'b0, 0, 0) c120131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120131));
	wire w320131;
	repeater #(1, 1'b0, 0, 0) c320131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320131));
	wire w930131;
	repeater #(1, 1'b1, 0, 0) c930131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w930131));
	wire w1270131;
	repeater #(1, 1'b1, 0, 0) c1270131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1270131));
	wire w1510131;

	wire w1520131;
	repeater #(1, 1'b0, 0, 0) c1520131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520131));
	wire w1590131;
	repeater #(2, 1'b1, 0, 0) c1590131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1590131));
	wire w1720131;
	assign outputs[73] = ();
	wire w1990131;
	repeater #(2, 1'b1, 0, 0) c1990131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990131));
	wire w2060131;
	repeater #(1, 1'b0, 0, 0) c2060131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060131));
	wire w2070131;

	wire w900133;
	torch #(1'b1) c900133 (.i_clk(tick), .i_in(), .o_out(w900133));
	wire w1060133;
	torch #(1'b1) c1060133 (.i_clk(tick), .i_in(), .o_out(w1060133));
	wire w1240133;
	torch #(1'b1) c1240133 (.i_clk(tick), .i_in(), .o_out(w1240133));
	wire w1400133;
	torch #(1'b1) c1400133 (.i_clk(tick), .i_in(), .o_out(w1400133));
	wire w980135;
	torch #(1'b1) c980135 (.i_clk(tick), .i_in(), .o_out(w980135));
	wire w1320135;
	torch #(1'b1) c1320135 (.i_clk(tick), .i_in(), .o_out(w1320135));
	wire w890136;
	repeater #(2, 1'b0, 0, 0) c890136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w890136));
	wire w1050136;
	repeater #(2, 1'b0, 0, 0) c1050136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1050136));
	wire w1230136;
	repeater #(2, 1'b0, 0, 0) c1230136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230136));
	wire w1390136;
	repeater #(2, 1'b0, 0, 0) c1390136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390136));
	wire w990137;
	repeater #(2, 1'b0, 0, 0) c990137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990137));
	wire w1330137;
	repeater #(2, 1'b0, 0, 0) c1330137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1330137));
	wire w80139;
	torch #(1'b1) c80139 (.i_clk(tick), .i_in(), .o_out(w80139));
	wire w120139;
	torch #(1'b1) c120139 (.i_clk(tick), .i_in(), .o_out(w120139));
	wire w160139;
	torch #(1'b1) c160139 (.i_clk(tick), .i_in(), .o_out(w160139));
	wire w200139;
	torch #(1'b1) c200139 (.i_clk(tick), .i_in(), .o_out(w200139));
	wire w240139;
	torch #(1'b1) c240139 (.i_clk(tick), .i_in(), .o_out(w240139));
	wire w280139;
	torch #(1'b1) c280139 (.i_clk(tick), .i_in(), .o_out(w280139));
	wire w320139;
	torch #(1'b1) c320139 (.i_clk(tick), .i_in(), .o_out(w320139));
	wire w60147;
	repeater #(1, 1'b0, 0, 0) c60147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60147));
	wire w120147;
	repeater #(1, 1'b0, 0, 0) c120147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120147));
	wire w320147;
	repeater #(1, 1'b0, 0, 0) c320147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320147));
	wire w1780153;

	wire w1790153;
	repeater #(1, 1'b0, 0, 0) c1790153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790153));
	wire w1800154;
	repeater #(1, 1'b0, 0, 0) c1800154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800154));
	wire w1830154;
	repeater #(2, 1'b0, 0, 0) c1830154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830154));
	wire w80155;
	torch #(1'b1) c80155 (.i_clk(tick), .i_in(), .o_out(w80155));
	wire w120155;
	torch #(1'b1) c120155 (.i_clk(tick), .i_in(), .o_out(w120155));
	wire w160155;
	torch #(1'b1) c160155 (.i_clk(tick), .i_in(), .o_out(w160155));
	wire w200155;
	torch #(1'b1) c200155 (.i_clk(tick), .i_in(), .o_out(w200155));
	wire w240155;
	torch #(1'b1) c240155 (.i_clk(tick), .i_in(), .o_out(w240155));
	wire w280155;
	torch #(1'b1) c280155 (.i_clk(tick), .i_in(), .o_out(w280155));
	wire w320155;
	torch #(1'b1) c320155 (.i_clk(tick), .i_in(), .o_out(w320155));
	wire w1750155;
	repeater #(1, 1'b0, 0, 0) c1750155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750155));
	wire w1880155;
	repeater #(2, 1'b0, 0, 0) c1880155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1880155));
	wire w1740156;
	assign outputs[74] = ();
	wire w1770156;

	wire w1860156;

	wire w1770157;

	wire w1860157;

	wire w1750158;
	repeater #(1, 1'b0, 0, 0) c1750158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750158));
	wire w1880158;
	repeater #(1, 1'b0, 0, 0) c1880158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1880158));
	wire w60163;
	repeater #(1, 1'b0, 0, 0) c60163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60163));
	wire w120163;
	repeater #(1, 1'b0, 0, 0) c120163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120163));
	wire w320163;
	repeater #(1, 1'b0, 0, 0) c320163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320163));
	wire w80171;
	torch #(1'b1) c80171 (.i_clk(tick), .i_in(), .o_out(w80171));
	wire w120171;
	torch #(1'b1) c120171 (.i_clk(tick), .i_in(), .o_out(w120171));
	wire w160171;
	torch #(1'b1) c160171 (.i_clk(tick), .i_in(), .o_out(w160171));
	wire w200171;
	torch #(1'b1) c200171 (.i_clk(tick), .i_in(), .o_out(w200171));
	wire w240171;
	torch #(1'b1) c240171 (.i_clk(tick), .i_in(), .o_out(w240171));
	wire w280171;
	torch #(1'b1) c280171 (.i_clk(tick), .i_in(), .o_out(w280171));
	wire w320171;
	torch #(1'b1) c320171 (.i_clk(tick), .i_in(), .o_out(w320171));
	wire w915;
	torch #(1'b1) c915 (.i_clk(tick), .i_in(), .o_out(w915));
	wire w1315;
	torch #(1'b1) c1315 (.i_clk(tick), .i_in(), .o_out(w1315));
	wire w1715;
	torch #(1'b1) c1715 (.i_clk(tick), .i_in(), .o_out(w1715));
	wire w2115;
	torch #(1'b1) c2115 (.i_clk(tick), .i_in(), .o_out(w2115));
	wire w2515;
	torch #(1'b1) c2515 (.i_clk(tick), .i_in(), .o_out(w2515));
	wire w2915;
	torch #(1'b1) c2915 (.i_clk(tick), .i_in(), .o_out(w2915));
	wire w3315;
	torch #(1'b1) c3315 (.i_clk(tick), .i_in(), .o_out(w3315));
	wire w919;
	torch #(1'b1) c919 (.i_clk(tick), .i_in(), .o_out(w919));
	wire w1319;
	torch #(1'b1) c1319 (.i_clk(tick), .i_in(), .o_out(w1319));
	wire w1719;
	torch #(1'b1) c1719 (.i_clk(tick), .i_in(), .o_out(w1719));
	wire w2119;
	torch #(1'b0) c2119 (.i_clk(tick), .i_in(), .o_out(w2119));
	wire w2519;
	torch #(1'b1) c2519 (.i_clk(tick), .i_in(), .o_out(w2519));
	wire w2919;
	torch #(1'b1) c2919 (.i_clk(tick), .i_in(), .o_out(w2919));
	wire w3319;
	torch #(1'b1) c3319 (.i_clk(tick), .i_in(), .o_out(w3319));
	wire w8117;
	torch #(1'b1) c8117 (.i_clk(tick), .i_in(), .o_out(w8117));
	wire w12117;
	torch #(1'b1) c12117 (.i_clk(tick), .i_in(), .o_out(w12117));
	wire w16117;
	torch #(1'b1) c16117 (.i_clk(tick), .i_in(), .o_out(w16117));
	wire w20117;
	torch #(1'b1) c20117 (.i_clk(tick), .i_in(), .o_out(w20117));
	wire w24117;
	torch #(1'b1) c24117 (.i_clk(tick), .i_in(), .o_out(w24117));
	wire w28117;
	torch #(1'b1) c28117 (.i_clk(tick), .i_in(), .o_out(w28117));
	wire w32117;
	torch #(1'b1) c32117 (.i_clk(tick), .i_in(), .o_out(w32117));
	wire w9150;
	repeater #(1, 1'b0, 0, 0) c9150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9150));
	wire w13150;
	repeater #(1, 1'b0, 0, 0) c13150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13150));
	wire w17150;
	repeater #(1, 1'b0, 0, 0) c17150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17150));
	wire w21150;
	repeater #(1, 1'b0, 0, 0) c21150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21150));
	wire w25150;
	repeater #(1, 1'b0, 0, 0) c25150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25150));
	wire w29150;
	repeater #(1, 1'b0, 0, 0) c29150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w29150));
	wire w33150;
	repeater #(1, 1'b0, 0, 0) c33150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33150));
	wire w9153;
	torch #(1'b1) c9153 (.i_clk(tick), .i_in(), .o_out(w9153));
	wire w13153;
	torch #(1'b1) c13153 (.i_clk(tick), .i_in(), .o_out(w13153));
	wire w17153;
	torch #(1'b1) c17153 (.i_clk(tick), .i_in(), .o_out(w17153));
	wire w21153;
	torch #(1'b1) c21153 (.i_clk(tick), .i_in(), .o_out(w21153));
	wire w25153;
	torch #(1'b1) c25153 (.i_clk(tick), .i_in(), .o_out(w25153));
	wire w29153;
	torch #(1'b1) c29153 (.i_clk(tick), .i_in(), .o_out(w29153));
	wire w33153;
	torch #(1'b1) c33153 (.i_clk(tick), .i_in(), .o_out(w33153));
	wire w20156;
	repeater #(1, 1'b1, 0, 0) c20156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20156));
	wire w22156;
	repeater #(1, 1'b1, 0, 0) c22156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22156));
	wire w24156;
	repeater #(1, 1'b1, 0, 0) c24156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24156));
	wire w26156;
	repeater #(1, 1'b1, 0, 0) c26156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26156));
	wire w28156;
	repeater #(1, 1'b1, 0, 0) c28156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28156));
	wire w30156;
	repeater #(1, 1'b1, 0, 0) c30156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30156));
	wire w32156;
	repeater #(1, 1'b1, 0, 0) c32156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32156));
	wire w34156;
	repeater #(1, 1'b1, 0, 0) c34156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34156));
	wire w18158;
	repeater #(1, 1'b1, 0, 0) c18158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18158));
	wire w16160;
	repeater #(1, 1'b1, 0, 0) c16160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16160));
	wire w14162;
	repeater #(1, 1'b1, 0, 0) c14162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14162));
	wire w12164;
	repeater #(1, 1'b1, 0, 0) c12164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12164));
	wire w10166;
	repeater #(1, 1'b1, 0, 0) c10166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10166));
	wire w8168;
	repeater #(1, 1'b1, 0, 0) c8168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8168));
	wire w106173;
	torch #(1'b1) c106173 (.i_clk(tick), .i_in(), .o_out(w106173));
	wire w140173;
	repeater #(1, 1'b1, 0, 0) c140173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140173));
	wire w174173;
	torch #(1'b1) c174173 (.i_clk(tick), .i_in(), .o_out(w174173));
	wire w0174;
	repeater #(1, 1'b1, 0, 0) c0174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0174));
	wire w104175;
	repeater #(1, 1'b0, 0, 0) c104175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104175));
	wire w138175;
	repeater #(1, 1'b0, 0, 0) c138175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138175));
	wire w172175;
	repeater #(1, 1'b1, 0, 0) c172175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172175));
	wire w206175;
	repeater #(1, 1'b1, 0, 0) c206175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206175));
	wire w34177;
	repeater #(1, 1'b1, 0, 0) c34177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34177));
	wire w102177;
	torch #(1'b1) c102177 (.i_clk(tick), .i_in(), .o_out(w102177));
	wire w136177;
	repeater #(1, 1'b1, 0, 0) c136177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136177));
	wire w170177;
	torch #(1'b1) c170177 (.i_clk(tick), .i_in(), .o_out(w170177));
	wire w204177;
	repeater #(1, 1'b1, 0, 0) c204177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204177));
	wire w32179;
	repeater #(1, 1'b1, 0, 0) c32179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32179));
	wire w100179;
	repeater #(1, 1'b1, 0, 0) c100179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100179));
	wire w134179;
	repeater #(1, 1'b1, 0, 0) c134179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134179));
	wire w168179;
	repeater #(1, 1'b1, 0, 0) c168179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168179));
	wire w202179;
	repeater #(1, 1'b1, 0, 0) c202179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202179));
	wire w30181;
	repeater #(1, 1'b1, 0, 0) c30181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30181));
	wire w98181;
	torch #(1'b1) c98181 (.i_clk(tick), .i_in(), .o_out(w98181));
	wire w132181;
	repeater #(1, 1'b1, 0, 0) c132181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132181));
	wire w166181;
	torch #(1'b1) c166181 (.i_clk(tick), .i_in(), .o_out(w166181));
	wire w200181;
	repeater #(1, 1'b1, 0, 0) c200181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200181));
	wire w28183;
	repeater #(1, 1'b1, 0, 0) c28183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w28183));
	wire w96183;
	repeater #(1, 1'b1, 0, 0) c96183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96183));
	wire w130183;
	repeater #(1, 1'b1, 0, 0) c130183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130183));
	wire w164183;
	repeater #(1, 1'b1, 0, 0) c164183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164183));
	wire w198183;
	repeater #(1, 1'b1, 0, 0) c198183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198183));
	wire w80184;
	repeater #(1, 1'b1, 0, 0) c80184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80184));
	wire w82184;
	torch #(1'b1) c82184 (.i_clk(tick), .i_in(), .o_out(w82184));
	wire w84184;
	repeater #(1, 1'b1, 0, 0) c84184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84184));
	wire w86184;
	torch #(1'b1) c86184 (.i_clk(tick), .i_in(), .o_out(w86184));
	wire w88184;
	repeater #(1, 1'b1, 0, 0) c88184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88184));
	wire w90184;
	torch #(1'b1) c90184 (.i_clk(tick), .i_in(), .o_out(w90184));
	wire w92184;
	repeater #(1, 1'b1, 0, 0) c92184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92184));
	wire w94184;
	torch #(1'b1) c94184 (.i_clk(tick), .i_in(), .o_out(w94184));
	wire w114184;
	repeater #(1, 1'b1, 0, 0) c114184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114184));
	wire w116184;
	repeater #(1, 1'b1, 0, 0) c116184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116184));
	wire w118184;
	repeater #(1, 1'b1, 0, 0) c118184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118184));
	wire w120184;
	repeater #(1, 1'b1, 0, 0) c120184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120184));
	wire w122184;
	repeater #(1, 1'b1, 0, 0) c122184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122184));
	wire w124184;
	repeater #(1, 1'b1, 0, 0) c124184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124184));
	wire w126184;
	repeater #(1, 1'b1, 0, 0) c126184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126184));
	wire w128184;
	repeater #(1, 1'b1, 0, 0) c128184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128184));
	wire w150184;
	torch #(1'b1) c150184 (.i_clk(tick), .i_in(), .o_out(w150184));
	wire w154184;
	torch #(1'b1) c154184 (.i_clk(tick), .i_in(), .o_out(w154184));
	wire w158184;
	torch #(1'b1) c158184 (.i_clk(tick), .i_in(), .o_out(w158184));
	wire w162184;
	torch #(1'b1) c162184 (.i_clk(tick), .i_in(), .o_out(w162184));
	wire w182184;
	repeater #(1, 1'b1, 0, 0) c182184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182184));
	wire w184184;
	repeater #(1, 1'b1, 0, 0) c184184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184184));
	wire w186184;
	repeater #(1, 1'b1, 0, 0) c186184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186184));
	wire w188184;
	repeater #(1, 1'b1, 0, 0) c188184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188184));
	wire w190184;
	repeater #(1, 1'b1, 0, 0) c190184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190184));
	wire w192184;
	repeater #(1, 1'b1, 0, 0) c192184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192184));
	wire w194184;
	repeater #(1, 1'b1, 0, 0) c194184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194184));
	wire w196184;
	repeater #(1, 1'b1, 0, 0) c196184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196184));
	wire w26185;
	repeater #(1, 1'b1, 0, 0) c26185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26185));
	wire w149185;
	repeater #(1, 1'b1, 0, 0) c149185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149185));
	wire w153185;
	repeater #(1, 1'b1, 0, 0) c153185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153185));
	wire w157185;
	repeater #(1, 1'b1, 0, 0) c157185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157185));
	wire w161185;
	repeater #(1, 1'b1, 0, 0) c161185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161185));
	wire w12186;
	repeater #(1, 1'b1, 0, 0) c12186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12186));
	wire w14186;
	repeater #(1, 1'b1, 0, 0) c14186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14186));
	wire w16186;
	repeater #(1, 1'b1, 0, 0) c16186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16186));
	wire w18186;
	repeater #(1, 1'b1, 0, 0) c18186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18186));
	wire w20186;
	repeater #(1, 1'b1, 0, 0) c20186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20186));
	wire w22186;
	repeater #(1, 1'b1, 0, 0) c22186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22186));
	wire w24186;
	repeater #(1, 1'b1, 0, 0) c24186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24186));
	wire w150187;
	torch #(1'b1) c150187 (.i_clk(tick), .i_in(), .o_out(w150187));
	wire w154187;
	torch #(1'b1) c154187 (.i_clk(tick), .i_in(), .o_out(w154187));
	wire w158187;
	torch #(1'b1) c158187 (.i_clk(tick), .i_in(), .o_out(w158187));
	wire w162187;
	torch #(1'b1) c162187 (.i_clk(tick), .i_in(), .o_out(w162187));
	wire w166187;
	torch #(1'b1) c166187 (.i_clk(tick), .i_in(), .o_out(w166187));
	wire w170187;
	torch #(1'b1) c170187 (.i_clk(tick), .i_in(), .o_out(w170187));
	wire w174187;
	torch #(1'b1) c174187 (.i_clk(tick), .i_in(), .o_out(w174187));
	wire w184187;
	torch #(1'b1) c184187 (.i_clk(tick), .i_in(), .o_out(w184187));
	wire w188187;
	torch #(1'b1) c188187 (.i_clk(tick), .i_in(), .o_out(w188187));
	wire w192187;
	torch #(1'b1) c192187 (.i_clk(tick), .i_in(), .o_out(w192187));
	wire w196187;
	torch #(1'b1) c196187 (.i_clk(tick), .i_in(), .o_out(w196187));
	wire w200187;
	torch #(1'b1) c200187 (.i_clk(tick), .i_in(), .o_out(w200187));
	wire w204187;
	torch #(1'b1) c204187 (.i_clk(tick), .i_in(), .o_out(w204187));
	wire w0188;
	torch #(1'b1) c0188 (.i_clk(tick), .i_in(), .o_out(w0188));
	wire w80188;
	repeater #(2, 1'b1, 0, 0) c80188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80188));
	wire w84188;
	repeater #(2, 1'b1, 0, 0) c84188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84188));
	wire w88188;
	repeater #(2, 1'b1, 0, 0) c88188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88188));
	wire w104188;
	repeater #(2, 1'b1, 0, 0) c104188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104188));
	wire w114188;
	repeater #(2, 1'b1, 0, 0) c114188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114188));
	wire w118188;
	repeater #(2, 1'b1, 0, 0) c118188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118188));
	wire w122188;
	repeater #(2, 1'b1, 0, 0) c122188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122188));
	wire w138188;
	repeater #(2, 1'b1, 0, 0) c138188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138188));
	wire w80190;
	torch #(1'b1) c80190 (.i_clk(tick), .i_in(), .o_out(w80190));
	wire w90190;
	repeater #(1, 1'b1, 0, 0) c90190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90190));
	wire w96190;
	torch #(1'b1) c96190 (.i_clk(tick), .i_in(), .o_out(w96190));
	wire w106190;
	repeater #(1, 1'b1, 0, 0) c106190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106190));
	wire w114190;
	torch #(1'b1) c114190 (.i_clk(tick), .i_in(), .o_out(w114190));
	wire w124190;
	repeater #(1, 1'b1, 0, 0) c124190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124190));
	wire w130190;
	torch #(1'b1) c130190 (.i_clk(tick), .i_in(), .o_out(w130190));
	wire w140190;
	repeater #(1, 1'b1, 0, 0) c140190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140190));
	wire w155191;
	torch #(1'b0) c155191 (.i_clk(tick), .i_in(), .o_out(w155191));
	wire w159191;
	torch #(1'b0) c159191 (.i_clk(tick), .i_in(), .o_out(w159191));
	wire w163191;
	torch #(1'b0) c163191 (.i_clk(tick), .i_in(), .o_out(w163191));
	wire w167191;
	torch #(1'b0) c167191 (.i_clk(tick), .i_in(), .o_out(w167191));
	wire w191191;
	torch #(1'b0) c191191 (.i_clk(tick), .i_in(), .o_out(w191191));
	wire w195191;
	torch #(1'b0) c195191 (.i_clk(tick), .i_in(), .o_out(w195191));
	wire w199191;
	torch #(1'b0) c199191 (.i_clk(tick), .i_in(), .o_out(w199191));
	wire w203191;
	torch #(1'b0) c203191 (.i_clk(tick), .i_in(), .o_out(w203191));
	wire w97193;
	repeater #(1, 1'b1, 0, 0) c97193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97193));
	wire w131193;
	repeater #(1, 1'b1, 0, 0) c131193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131193));
	wire w90194;
	repeater #(1, 1'b1, 0, 0) c90194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90194));
	wire w103194;

	wire w106194;
	repeater #(1, 1'b1, 0, 0) c106194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106194));
	wire w124194;
	repeater #(1, 1'b1, 0, 0) c124194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124194));
	wire w137194;

	wire w140194;
	repeater #(1, 1'b1, 0, 0) c140194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140194));
	wire w79195;

	wire w95195;

	wire w113195;

	wire w129195;

	wire w10196;
	repeater #(1, 1'b1, 0, 0) c10196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10196));
	wire w14196;
	repeater #(1, 1'b1, 0, 0) c14196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14196));
	wire w18196;
	repeater #(1, 1'b1, 0, 0) c18196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18196));
	wire w22196;
	repeater #(1, 1'b1, 0, 0) c22196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22196));
	wire w26196;
	repeater #(1, 1'b1, 0, 0) c26196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26196));
	wire w30196;
	repeater #(1, 1'b1, 0, 0) c30196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30196));
	wire w34196;
	repeater #(1, 1'b1, 0, 0) c34196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34196));
	wire w103196;

	wire w137196;

	wire w89197;

	wire w90197;

	wire w100197;

	wire w105197;

	wire w106197;

	wire w123197;

	wire w124197;

	wire w134197;

	wire w139197;

	wire w140197;

	wire w82199;

	wire w98199;

	wire w116199;

	wire w132199;

	wire w121100;

	wire w371100;
	repeater #(2, 1'b0, 0, 0) c371100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w371100));
	wire w881100;

	wire w891100;

	wire w1041100;

	wire w1051100;

	wire w1221100;

	wire w1231100;

	wire w1381100;

	wire w1391100;

	wire w321101;

	wire w981101;

	wire w1021101;

	wire w1321101;

	wire w1361101;

	wire w71102;
	repeater #(1, 1'b0, 0, 0) c71102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71102));
	wire w161105;
	torch #(1'b1) c161105 (.i_clk(tick), .i_in(), .o_out(w161105));
	wire w201105;
	torch #(1'b1) c201105 (.i_clk(tick), .i_in(), .o_out(w201105));
	wire w241105;
	torch #(1'b1) c241105 (.i_clk(tick), .i_in(), .o_out(w241105));
	wire w281105;
	torch #(1'b1) c281105 (.i_clk(tick), .i_in(), .o_out(w281105));
	wire w791105;

	wire w801105;

	wire w831105;

	wire w841105;

	wire w871105;

	wire w881105;

	wire w911105;

	wire w921105;

	wire w951105;

	wire w961105;

	wire w991105;

	wire w1001105;

	wire w1031105;

	wire w1041105;

	wire w1131105;

	wire w1141105;

	wire w1171105;

	wire w1181105;

	wire w1211105;

	wire w1221105;

	wire w1251105;

	wire w1261105;

	wire w1291105;

	wire w1301105;

	wire w1331105;

	wire w1341105;

	wire w1371105;

	wire w1381105;

	wire w801107;

	wire w841107;

	wire w881107;

	wire w921107;

	wire w961107;

	wire w1001107;

	wire w1041107;

	wire w1141107;

	wire w1181107;

	wire w1221107;

	wire w1261107;

	wire w1301107;

	wire w1341107;

	wire w1381107;

	wire w91109;
	torch #(1'b0) c91109 (.i_clk(tick), .i_in(), .o_out(w91109));
	wire w131109;
	torch #(1'b0) c131109 (.i_clk(tick), .i_in(), .o_out(w131109));
	wire w171109;
	torch #(1'b0) c171109 (.i_clk(tick), .i_in(), .o_out(w171109));
	wire w211109;
	torch #(1'b0) c211109 (.i_clk(tick), .i_in(), .o_out(w211109));
	wire w251109;
	torch #(1'b0) c251109 (.i_clk(tick), .i_in(), .o_out(w251109));
	wire w291109;
	torch #(1'b0) c291109 (.i_clk(tick), .i_in(), .o_out(w291109));
	wire w331109;
	torch #(1'b0) c331109 (.i_clk(tick), .i_in(), .o_out(w331109));
	wire w781110;

	wire w821110;

	wire w861110;

	wire w901110;

	wire w1121110;

	wire w1161110;

	wire w1201110;

	wire w1241110;

	wire w101111;
	torch #(1'b1) c101111 (.i_clk(tick), .i_in(), .o_out(w101111));
	wire w141111;
	torch #(1'b1) c141111 (.i_clk(tick), .i_in(), .o_out(w141111));
	wire w181111;
	torch #(1'b1) c181111 (.i_clk(tick), .i_in(), .o_out(w181111));
	wire w221111;
	torch #(1'b1) c221111 (.i_clk(tick), .i_in(), .o_out(w221111));
	wire w261111;
	torch #(1'b1) c261111 (.i_clk(tick), .i_in(), .o_out(w261111));
	wire w301111;
	torch #(1'b1) c301111 (.i_clk(tick), .i_in(), .o_out(w301111));
	wire w341111;
	torch #(1'b1) c341111 (.i_clk(tick), .i_in(), .o_out(w341111));
	wire w901112;

	wire w1241112;

	wire w881113;
	repeater #(1, 1'b1, 0, 0) c881113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w881113));
	wire w1221113;
	repeater #(1, 1'b1, 0, 0) c1221113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221113));
	wire w791114;
	repeater #(1, 1'b1, 0, 0) c791114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791114));
	wire w821114;

	wire w951114;
	repeater #(1, 1'b1, 0, 0) c951114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951114));
	wire w1131114;
	repeater #(1, 1'b1, 0, 0) c1131114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1131114));
	wire w1161114;

	wire w1291114;
	repeater #(1, 1'b1, 0, 0) c1291114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1291114));
	wire w901115;

	wire w1241115;

	wire w121116;

	wire w371116;
	repeater #(2, 1'b0, 0, 0) c371116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w371116));
	wire w821116;

	wire w1161116;

	wire w321117;

	wire w791117;

	wire w801117;

	wire w851117;

	wire w931117;

	wire w951117;

	wire w1131117;

	wire w1141117;

	wire w1191117;

	wire w1271117;

	wire w1291117;

	wire w71118;
	repeater #(1, 1'b0, 0, 0) c71118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71118));
	wire w871119;

	wire w881119;

	wire w1211119;

	wire w1221119;

	wire w1701119;
	repeater #(1, 1'b1, 0, 0) c1701119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701119));
	wire w1881119;
	repeater #(1, 1'b1, 0, 0) c1881119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1881119));
	wire w161121;
	torch #(1'b1) c161121 (.i_clk(tick), .i_in(), .o_out(w161121));
	wire w201121;
	torch #(1'b1) c201121 (.i_clk(tick), .i_in(), .o_out(w201121));
	wire w241121;
	torch #(1'b1) c241121 (.i_clk(tick), .i_in(), .o_out(w241121));
	wire w281121;
	torch #(1'b1) c281121 (.i_clk(tick), .i_in(), .o_out(w281121));
	wire w791121;

	wire w801121;

	wire w931121;

	wire w951121;

	wire w961121;

	wire w1131121;

	wire w1141121;

	wire w1271121;

	wire w1291121;

	wire w1301121;

	wire w1771122;
	repeater #(1, 1'b1, 0, 0) c1771122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1771122));
	wire w901123;
	torch #(1'b1) c901123 (.i_clk(tick), .i_in(), .o_out(w901123));
	wire w911123;

	wire w1241123;
	torch #(1'b1) c1241123 (.i_clk(tick), .i_in(), .o_out(w1241123));
	wire w1251123;

	wire w911124;

	wire w931124;

	wire w1251124;

	wire w1271124;

	wire w1491124;
	repeater #(1, 1'b1, 0, 0) c1491124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1491124));
	wire w1811124;

	wire w11125;
	repeater #(1, 1'b0, 0, 0) c11125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11125));
	wire w91125;
	torch #(1'b0) c91125 (.i_clk(tick), .i_in(), .o_out(w91125));
	wire w131125;
	torch #(1'b0) c131125 (.i_clk(tick), .i_in(), .o_out(w131125));
	wire w171125;
	torch #(1'b0) c171125 (.i_clk(tick), .i_in(), .o_out(w171125));
	wire w211125;
	torch #(1'b0) c211125 (.i_clk(tick), .i_in(), .o_out(w211125));
	wire w251125;
	torch #(1'b0) c251125 (.i_clk(tick), .i_in(), .o_out(w251125));
	wire w291125;
	torch #(1'b0) c291125 (.i_clk(tick), .i_in(), .o_out(w291125));
	wire w331125;
	torch #(1'b0) c331125 (.i_clk(tick), .i_in(), .o_out(w331125));
	wire w1531125;
	repeater #(1, 1'b1, 0, 0) c1531125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1531125));
	wire w1781125;

	wire w2051125;
	repeater #(1, 1'b0, 0, 0) c2051125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2051125));
	wire w931126;

	wire w941126;

	wire w951126;

	wire w1271126;

	wire w1281126;

	wire w1291126;

	wire w1591126;

	wire w1631126;
	repeater #(1, 1'b0, 0, 0) c1631126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1631126));
	wire w1771126;

	wire w1791126;
	repeater #(2, 1'b1, 0, 0) c1791126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1791126));
	wire w1821126;
	repeater #(2, 1'b1, 0, 0) c1821126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821126));
	wire w1951126;
	repeater #(1, 1'b0, 0, 0) c1951126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1951126));
	wire w1991126;

	wire w101127;
	torch #(1'b1) c101127 (.i_clk(tick), .i_in(), .o_out(w101127));
	wire w141127;
	torch #(1'b1) c141127 (.i_clk(tick), .i_in(), .o_out(w141127));
	wire w181127;
	torch #(1'b1) c181127 (.i_clk(tick), .i_in(), .o_out(w181127));
	wire w221127;
	torch #(1'b1) c221127 (.i_clk(tick), .i_in(), .o_out(w221127));
	wire w261127;
	torch #(1'b1) c261127 (.i_clk(tick), .i_in(), .o_out(w261127));
	wire w301127;
	torch #(1'b1) c301127 (.i_clk(tick), .i_in(), .o_out(w301127));
	wire w341127;
	torch #(1'b1) c341127 (.i_clk(tick), .i_in(), .o_out(w341127));
	wire w881127;

	wire w891127;

	wire w951127;

	wire w1041127;

	wire w1051127;

	wire w1221127;

	wire w1231127;

	wire w1291127;

	wire w1381127;

	wire w1391127;

	wire w1601127;

	wire w1661127;
	repeater #(2, 1'b0, 0, 0) c1661127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661127));
	wire w1691127;
	repeater #(2, 1'b0, 0, 0) c1691127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1691127));
	wire w1711127;

	wire w1871127;

	wire w1891127;
	repeater #(2, 1'b0, 0, 0) c1891127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1891127));
	wire w1921127;
	repeater #(2, 1'b0, 0, 0) c1921127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1921127));
	wire w1981127;

	wire w1591128;
	repeater #(2, 1'b1, 0, 0) c1591128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591128));
	wire w1701128;

	wire w1881128;

	wire w1991128;
	repeater #(2, 1'b0, 0, 0) c1991128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991128));
	wire w931129;
	repeater #(1, 1'b0, 0, 0) c931129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w931129));
	wire w951129;
	torch #(1'b0) c951129 (.i_clk(tick), .i_in(), .o_out(w951129));
	wire w1011129;
	torch #(1'b0) c1011129 (.i_clk(tick), .i_in(), .o_out(w1011129));
	wire w1271129;
	repeater #(1, 1'b0, 0, 0) c1271129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271129));
	wire w1291129;
	torch #(1'b0) c1291129 (.i_clk(tick), .i_in(), .o_out(w1291129));
	wire w1351129;
	torch #(1'b0) c1351129 (.i_clk(tick), .i_in(), .o_out(w1351129));
	wire w1531129;

	wire w1541129;

	wire w1671129;

	wire w1911129;

	wire w2041129;

	wire w2051129;

	wire w1521130;

	wire w1611130;

	wire w1971130;

	wire w2061130;

	wire w971131;
	repeater #(1, 1'b1, 0, 0) c971131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w971131));
	wire w1311131;
	repeater #(1, 1'b1, 0, 0) c1311131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1311131));
	wire w1851131;
	assign outputs[75] = ();
	wire w121132;

	wire w371132;
	repeater #(2, 1'b0, 0, 0) c371132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w371132));
	wire w321133;

	wire w941133;
	torch #(1'b1) c941133 (.i_clk(tick), .i_in(), .o_out(w941133));
	wire w1281133;
	torch #(1'b1) c1281133 (.i_clk(tick), .i_in(), .o_out(w1281133));
	wire w71134;
	repeater #(1, 1'b0, 0, 0) c71134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71134));
	wire w1021135;
	torch #(1'b1) c1021135 (.i_clk(tick), .i_in(), .o_out(w1021135));
	wire w1361135;
	torch #(1'b1) c1361135 (.i_clk(tick), .i_in(), .o_out(w1361135));
	wire w7700;
	repeater #(2, 1'b0, 0, 0) c7700 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7700));
	wire w11100;
	repeater #(2, 1'b0, 0, 0) c11100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11100));
	wire w001;
	torch #(1'b1) c001 (.i_clk(tick), .i_in(), .o_out(w001));
	wire w401;
	torch #(1'b1) c401 (.i_clk(tick), .i_in(), .o_out(w401));
	wire w801;
	torch #(1'b1) c801 (.i_clk(tick), .i_in(), .o_out(w801));
	wire w1201;
	torch #(1'b1) c1201 (.i_clk(tick), .i_in(), .o_out(w1201));
	wire w8701;
	repeater #(2, 1'b0, 0, 0) c8701 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8701));
	wire w12101;
	repeater #(2, 1'b0, 0, 0) c12101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12101));
	wire w20104;
	torch #(1'b0) c20104 (.i_clk(tick), .i_in(), .o_out(w20104));
	wire w20504;
	torch #(1'b0) c20504 (.i_clk(tick), .i_in(), .o_out(w20504));
	wire w105;
	torch #(1'b0) c105 (.i_clk(tick), .i_in(), .o_out(w105));
	wire w505;
	torch #(1'b0) c505 (.i_clk(tick), .i_in(), .o_out(w505));
	wire w905;
	torch #(1'b0) c905 (.i_clk(tick), .i_in(), .o_out(w905));
	wire w1305;
	torch #(1'b0) c1305 (.i_clk(tick), .i_in(), .o_out(w1305));
	wire w1705;
	torch #(1'b0) c1705 (.i_clk(tick), .i_in(), .o_out(w1705));
	wire w20206;
	torch #(1'b1) c20206 (.i_clk(tick), .i_in(), .o_out(w20206));
	wire w20606;
	torch #(1'b1) c20606 (.i_clk(tick), .i_in(), .o_out(w20606));
	wire w207;
	torch #(1'b1) c207 (.i_clk(tick), .i_in(), .o_out(w207));
	wire w607;
	torch #(1'b1) c607 (.i_clk(tick), .i_in(), .o_out(w607));
	wire w1007;
	torch #(1'b1) c1007 (.i_clk(tick), .i_in(), .o_out(w1007));
	wire w1407;
	torch #(1'b1) c1407 (.i_clk(tick), .i_in(), .o_out(w1407));
	wire w1807;
	torch #(1'b1) c1807 (.i_clk(tick), .i_in(), .o_out(w1807));
	wire w97010;
	repeater #(1, 1'b0, 0, 0) c97010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97010));
	wire w84011;
	repeater #(1, 1'b0, 0, 0) c84011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84011));
	wire w104011;
	repeater #(2, 1'b0, 0, 0) c104011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104011));
	wire w204011;

	wire w21012;
	repeater #(2, 1'b0, 0, 0) c21012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21012));
	wire w16013;

	wire w199013;
	repeater #(1, 1'b0, 0, 0) c199013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199013));
	wire w0017;
	torch #(1'b1) c0017 (.i_clk(tick), .i_in(), .o_out(w0017));
	wire w4017;
	torch #(1'b1) c4017 (.i_clk(tick), .i_in(), .o_out(w4017));
	wire w8017;
	torch #(1'b1) c8017 (.i_clk(tick), .i_in(), .o_out(w8017));
	wire w12017;
	torch #(1'b1) c12017 (.i_clk(tick), .i_in(), .o_out(w12017));
	wire w156017;

	wire w174017;

	wire w201020;
	torch #(1'b0) c201020 (.i_clk(tick), .i_in(), .o_out(w201020));
	wire w205020;
	torch #(1'b0) c205020 (.i_clk(tick), .i_in(), .o_out(w205020));
	wire w1021;
	torch #(1'b0) c1021 (.i_clk(tick), .i_in(), .o_out(w1021));
	wire w5021;
	torch #(1'b0) c5021 (.i_clk(tick), .i_in(), .o_out(w5021));
	wire w9021;
	torch #(1'b0) c9021 (.i_clk(tick), .i_in(), .o_out(w9021));
	wire w13021;
	torch #(1'b0) c13021 (.i_clk(tick), .i_in(), .o_out(w13021));
	wire w17021;
	torch #(1'b0) c17021 (.i_clk(tick), .i_in(), .o_out(w17021));
	wire w202022;
	torch #(1'b1) c202022 (.i_clk(tick), .i_in(), .o_out(w202022));
	wire w206022;
	torch #(1'b1) c206022 (.i_clk(tick), .i_in(), .o_out(w206022));
	wire w2023;
	torch #(1'b1) c2023 (.i_clk(tick), .i_in(), .o_out(w2023));
	wire w6023;
	torch #(1'b1) c6023 (.i_clk(tick), .i_in(), .o_out(w6023));
	wire w10023;
	torch #(1'b1) c10023 (.i_clk(tick), .i_in(), .o_out(w10023));
	wire w14023;
	torch #(1'b1) c14023 (.i_clk(tick), .i_in(), .o_out(w14023));
	wire w18023;
	torch #(1'b1) c18023 (.i_clk(tick), .i_in(), .o_out(w18023));
	wire w204027;

	wire w21028;
	repeater #(2, 1'b0, 0, 0) c21028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21028));
	wire w16029;

	wire w199029;
	repeater #(1, 1'b0, 0, 0) c199029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199029));
	wire w0033;
	torch #(1'b1) c0033 (.i_clk(tick), .i_in(), .o_out(w0033));
	wire w4033;
	torch #(1'b1) c4033 (.i_clk(tick), .i_in(), .o_out(w4033));
	wire w8033;
	torch #(1'b1) c8033 (.i_clk(tick), .i_in(), .o_out(w8033));
	wire w12033;
	torch #(1'b1) c12033 (.i_clk(tick), .i_in(), .o_out(w12033));
	wire w201036;
	torch #(1'b0) c201036 (.i_clk(tick), .i_in(), .o_out(w201036));
	wire w205036;
	torch #(1'b0) c205036 (.i_clk(tick), .i_in(), .o_out(w205036));
	wire w1037;
	torch #(1'b0) c1037 (.i_clk(tick), .i_in(), .o_out(w1037));
	wire w5037;
	torch #(1'b0) c5037 (.i_clk(tick), .i_in(), .o_out(w5037));
	wire w9037;
	torch #(1'b0) c9037 (.i_clk(tick), .i_in(), .o_out(w9037));
	wire w13037;
	torch #(1'b0) c13037 (.i_clk(tick), .i_in(), .o_out(w13037));
	wire w17037;
	torch #(1'b0) c17037 (.i_clk(tick), .i_in(), .o_out(w17037));
	wire w202038;
	torch #(1'b1) c202038 (.i_clk(tick), .i_in(), .o_out(w202038));
	wire w206038;
	torch #(1'b1) c206038 (.i_clk(tick), .i_in(), .o_out(w206038));
	wire w2039;
	torch #(1'b1) c2039 (.i_clk(tick), .i_in(), .o_out(w2039));
	wire w6039;
	torch #(1'b1) c6039 (.i_clk(tick), .i_in(), .o_out(w6039));
	wire w10039;
	torch #(1'b1) c10039 (.i_clk(tick), .i_in(), .o_out(w10039));
	wire w14039;
	torch #(1'b1) c14039 (.i_clk(tick), .i_in(), .o_out(w14039));
	wire w18039;
	torch #(1'b1) c18039 (.i_clk(tick), .i_in(), .o_out(w18039));
	wire w199050;
	repeater #(2, 1'b0, 0, 0) c199050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199050));
	wire w203050;
	repeater #(2, 1'b0, 0, 0) c203050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203050));
	wire w207050;
	repeater #(2, 1'b0, 0, 0) c207050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207050));
	wire w3051;
	repeater #(2, 1'b0, 0, 0) c3051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3051));
	wire w7051;
	repeater #(2, 1'b0, 0, 0) c7051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7051));
	wire w11051;
	repeater #(2, 1'b0, 0, 0) c11051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11051));
	wire w15051;
	repeater #(2, 1'b0, 0, 0) c15051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15051));
	wire w200052;

	wire w204052;

	wire w0053;

	wire w4053;

	wire w8053;

	wire w12053;

	wire w16053;

	wire w200053;

	wire w204053;

	wire w0054;

	wire w4054;

	wire w8054;

	wire w12054;

	wire w16054;

	wire w199056;
	repeater #(1, 1'b1, 0, 0) c199056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199056));
	wire w203056;
	repeater #(1, 1'b1, 0, 0) c203056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203056));
	wire w207056;
	repeater #(1, 1'b1, 0, 0) c207056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207056));
	wire w3057;
	repeater #(1, 1'b0, 0, 0) c3057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3057));
	wire w7057;
	repeater #(1, 1'b1, 0, 0) c7057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7057));
	wire w11057;
	repeater #(1, 1'b1, 0, 0) c11057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11057));
	wire w15057;
	repeater #(1, 1'b1, 0, 0) c15057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15057));
	wire w201057;

	wire w205057;

	wire w1058;

	wire w5058;

	wire w9058;

	wire w13058;

	wire w17058;

	wire w200058;

	wire w204058;

	wire w0059;

	wire w4059;

	wire w8059;

	wire w12059;

	wire w16059;

	wire w202060;
	torch #(1'b0) c202060 (.i_clk(tick), .i_in(), .o_out(w202060));
	wire w206060;
	torch #(1'b0) c206060 (.i_clk(tick), .i_in(), .o_out(w206060));
	wire w2061;
	torch #(1'b0) c2061 (.i_clk(tick), .i_in(), .o_out(w2061));
	wire w6061;
	torch #(1'b1) c6061 (.i_clk(tick), .i_in(), .o_out(w6061));
	wire w10061;
	torch #(1'b0) c10061 (.i_clk(tick), .i_in(), .o_out(w10061));
	wire w14061;
	torch #(1'b0) c14061 (.i_clk(tick), .i_in(), .o_out(w14061));
	wire w18061;
	torch #(1'b0) c18061 (.i_clk(tick), .i_in(), .o_out(w18061));
	wire w24063;
	repeater #(1, 1'b1, 0, 0) c24063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24063));
	wire w90099;

	wire w123099;

	wire w124099;

	wire w157099;

	wire w158099;

	wire w191099;

	wire w192099;

	wire w170100;

	wire w910100;
	repeater #(1, 1'b1, 0, 0) c910100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w910100));
	wire w1250100;
	repeater #(1, 1'b1, 0, 0) c1250100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1250100));
	wire w1590100;
	repeater #(1, 1'b1, 0, 0) c1590100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1590100));
	wire w1930100;
	repeater #(1, 1'b1, 0, 0) c1930100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1930100));
	wire w880101;

	wire w1210101;

	wire w1220101;

	wire w1550101;

	wire w1560101;

	wire w1890101;

	wire w1900101;

	wire w150102;

	wire w180102;
	repeater #(1, 1'b1, 0, 0) c180102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180102));
	wire w890102;
	repeater #(1, 1'b0, 0, 0) c890102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w890102));
	wire w1230102;
	repeater #(1, 1'b0, 0, 0) c1230102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230102));
	wire w1570102;
	repeater #(1, 1'b1, 0, 0) c1570102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570102));
	wire w1910102;
	repeater #(1, 1'b1, 0, 0) c1910102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910102));
	wire w170103;

	wire w860103;

	wire w1190103;

	wire w1200103;

	wire w1530103;

	wire w1540103;

	wire w1870103;

	wire w1880103;

	wire w130104;

	wire w160104;
	repeater #(1, 1'b1, 0, 0) c160104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160104));
	wire w870104;
	repeater #(1, 1'b1, 0, 0) c870104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w870104));
	wire w1210104;
	repeater #(1, 1'b1, 0, 0) c1210104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1210104));
	wire w1550104;
	repeater #(1, 1'b1, 0, 0) c1550104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550104));
	wire w1890104;
	repeater #(1, 1'b1, 0, 0) c1890104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1890104));
	wire w150105;

	wire w840105;

	wire w1170105;

	wire w1180105;

	wire w1510105;

	wire w1520105;

	wire w1850105;

	wire w1860105;

	wire w110106;

	wire w140106;
	repeater #(1, 1'b1, 0, 0) c140106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140106));
	wire w850106;
	repeater #(1, 1'b1, 0, 0) c850106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w850106));
	wire w1190106;
	repeater #(1, 1'b1, 0, 0) c1190106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190106));
	wire w1530106;
	repeater #(1, 1'b1, 0, 0) c1530106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1530106));
	wire w1870106;
	repeater #(1, 1'b1, 0, 0) c1870106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870106));
	wire w130107;

	wire w820107;

	wire w1150107;

	wire w1160107;

	wire w1490107;

	wire w1500107;

	wire w1830107;

	wire w1840107;

	wire w90108;

	wire w120108;
	repeater #(1, 1'b1, 0, 0) c120108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120108));
	wire w830108;
	repeater #(1, 1'b1, 0, 0) c830108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w830108));
	wire w1170108;
	repeater #(1, 1'b1, 0, 0) c1170108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1170108));
	wire w1510108;
	repeater #(1, 1'b1, 0, 0) c1510108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510108));
	wire w1850108;
	repeater #(1, 1'b1, 0, 0) c1850108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850108));
	wire w110109;

	wire w800109;

	wire w1130109;

	wire w1140109;

	wire w1470109;

	wire w1480109;

	wire w1810109;

	wire w1820109;

	wire w70110;

	wire w100110;
	repeater #(1, 1'b1, 0, 0) c100110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100110));
	wire w810110;
	repeater #(1, 1'b1, 0, 0) c810110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w810110));
	wire w1150110;
	repeater #(1, 1'b1, 0, 0) c1150110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1150110));
	wire w1490110;
	repeater #(1, 1'b1, 0, 0) c1490110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490110));
	wire w1830110;
	repeater #(1, 1'b1, 0, 0) c1830110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830110));
	wire w90111;

	wire w780111;

	wire w1110111;

	wire w1120111;

	wire w1450111;

	wire w1460111;

	wire w1790111;

	wire w1800111;

	wire w50112;

	wire w80112;
	repeater #(1, 1'b1, 0, 0) c80112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80112));
	wire w790112;
	repeater #(1, 1'b1, 0, 0) c790112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w790112));
	wire w1130112;
	repeater #(1, 1'b1, 0, 0) c1130112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1130112));
	wire w1470112;
	repeater #(1, 1'b1, 0, 0) c1470112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470112));
	wire w1810112;
	repeater #(1, 1'b1, 0, 0) c1810112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810112));
	wire w70113;

	wire w760113;

	wire w1090113;

	wire w1100113;

	wire w1430113;

	wire w1440113;

	wire w1770113;

	wire w1780113;

	wire w30114;

	wire w60114;
	repeater #(1, 1'b1, 0, 0) c60114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60114));
	wire w770114;
	repeater #(1, 1'b1, 0, 0) c770114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w770114));
	wire w1110114;
	repeater #(1, 1'b1, 0, 0) c1110114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110114));
	wire w1450114;
	repeater #(1, 1'b1, 0, 0) c1450114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450114));
	wire w1790114;
	repeater #(1, 1'b1, 0, 0) c1790114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790114));
	wire w50115;

	wire w740115;

	wire w1070115;

	wire w1080115;

	wire w1410115;

	wire w1420115;

	wire w1750115;

	wire w1760115;

	wire w10116;

	wire w40116;
	repeater #(1, 1'b1, 0, 0) c40116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40116));
	wire w750116;
	repeater #(1, 1'b1, 0, 0) c750116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w750116));
	wire w1090116;
	repeater #(1, 1'b1, 0, 0) c1090116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1090116));
	wire w1430116;
	repeater #(1, 1'b1, 0, 0) c1430116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1430116));
	wire w1770116;
	repeater #(1, 1'b1, 0, 0) c1770116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770116));
	wire w30117;

	wire w720117;

	wire w1050117;

	wire w1060117;

	wire w1390117;

	wire w1400117;

	wire w1730117;

	wire w1740117;

	wire w2070117;

	wire w20118;
	repeater #(1, 1'b1, 0, 0) c20118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20118));
	wire w730118;
	repeater #(1, 1'b1, 0, 0) c730118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w730118));
	wire w1070118;
	repeater #(1, 1'b1, 0, 0) c1070118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1070118));
	wire w1410118;
	repeater #(1, 1'b1, 0, 0) c1410118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1410118));
	wire w1750118;
	repeater #(1, 1'b1, 0, 0) c1750118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750118));
	wire w10119;

	wire w700119;

	wire w1030119;

	wire w1040119;

	wire w1370119;

	wire w1380119;

	wire w1710119;

	wire w1720119;

	wire w2050119;

	wire w00120;
	repeater #(1, 1'b1, 0, 0) c00120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w00120));
	wire w710120;
	repeater #(1, 1'b1, 0, 0) c710120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w710120));
	wire w1050120;
	repeater #(1, 1'b1, 0, 0) c1050120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1050120));
	wire w1390120;
	repeater #(1, 1'b1, 0, 0) c1390120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390120));
	wire w1730120;
	repeater #(1, 1'b1, 0, 0) c1730120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1730120));
	wire w2070120;

	wire w680121;

	wire w1010121;

	wire w1020121;

	wire w1350121;

	wire w1360121;

	wire w1690121;

	wire w1700121;

	wire w2030121;

	wire w2060121;
	repeater #(1, 1'b1, 0, 0) c2060121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060121));
	wire w690122;
	repeater #(1, 1'b1, 0, 0) c690122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w690122));
	wire w1030122;
	repeater #(1, 1'b1, 0, 0) c1030122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1030122));
	wire w1370122;
	repeater #(1, 1'b1, 0, 0) c1370122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370122));
	wire w1710122;
	repeater #(1, 1'b1, 0, 0) c1710122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710122));
	wire w2050122;

	wire w660123;

	wire w990123;

	wire w1000123;

	wire w1330123;

	wire w1340123;

	wire w1670123;

	wire w1680123;

	wire w2010123;

	wire w2040123;
	repeater #(1, 1'b1, 0, 0) c2040123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2040123));
	wire w670124;
	repeater #(1, 1'b1, 0, 0) c670124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w670124));
	wire w1010124;
	repeater #(1, 1'b1, 0, 0) c1010124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010124));
	wire w1350124;
	repeater #(1, 1'b1, 0, 0) c1350124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350124));
	wire w1690124;
	repeater #(1, 1'b1, 0, 0) c1690124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1690124));
	wire w2030124;

	wire w970125;

	wire w1310125;

	wire w1650125;

	wire w1990125;

	wire w2020125;
	repeater #(1, 1'b1, 0, 0) c2020125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020125));
	wire w650126;
	repeater #(1, 1'b1, 0, 0) c650126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650126));
	wire w990126;
	repeater #(1, 1'b1, 0, 0) c990126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w990126));
	wire w1330126;
	repeater #(1, 1'b1, 0, 0) c1330126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1330126));
	wire w1670126;
	repeater #(1, 1'b1, 0, 0) c1670126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1670126));
	wire w2010126;

	wire w2000127;
	repeater #(2, 1'b1, 0, 0) c2000127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2000127));
	wire w2020128;
	repeater #(1, 1'b1, 0, 0) c2020128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020128));
	wire w840131;
	repeater #(2, 1'b1, 0, 0) c840131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840131));
	wire w1180131;
	repeater #(2, 1'b1, 0, 0) c1180131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1180131));
	wire w2010131;
	torch #(1'b1) c2010131 (.i_clk(tick), .i_in(), .o_out(w2010131));
	wire w2050131;
	torch #(1'b1) c2050131 (.i_clk(tick), .i_in(), .o_out(w2050131));
	wire w10132;
	torch #(1'b1) c10132 (.i_clk(tick), .i_in(), .o_out(w10132));
	wire w50132;
	torch #(1'b1) c50132 (.i_clk(tick), .i_in(), .o_out(w50132));
	wire w90132;
	torch #(1'b1) c90132 (.i_clk(tick), .i_in(), .o_out(w90132));
	wire w130132;
	torch #(1'b1) c130132 (.i_clk(tick), .i_in(), .o_out(w130132));
	wire w170132;
	torch #(1'b1) c170132 (.i_clk(tick), .i_in(), .o_out(w170132));
	wire w700133;
	repeater #(1, 1'b1, 0, 0) c700133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w700133));
	wire w760133;
	torch #(1'b1) c760133 (.i_clk(tick), .i_in(), .o_out(w760133));
	wire w860133;
	repeater #(1, 1'b1, 0, 0) c860133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w860133));
	wire w1040133;
	repeater #(1, 1'b1, 0, 0) c1040133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1040133));
	wire w1100133;
	torch #(1'b1) c1100133 (.i_clk(tick), .i_in(), .o_out(w1100133));
	wire w1200133;
	repeater #(1, 1'b1, 0, 0) c1200133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1200133));
	wire w2020134;
	repeater #(1, 1'b1, 0, 0) c2020134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020134));
	wire w2060134;
	repeater #(1, 1'b1, 0, 0) c2060134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060134));
	wire w20135;
	repeater #(1, 1'b1, 0, 0) c20135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20135));
	wire w60135;
	repeater #(1, 1'b1, 0, 0) c60135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60135));
	wire w100135;
	repeater #(1, 1'b1, 0, 0) c100135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100135));
	wire w140135;
	repeater #(1, 1'b1, 0, 0) c140135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140135));
	wire w180135;
	repeater #(1, 1'b1, 0, 0) c180135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180135));
	wire w2010135;
	torch #(1'b1) c2010135 (.i_clk(tick), .i_in(), .o_out(w2010135));
	wire w2050135;
	torch #(1'b1) c2050135 (.i_clk(tick), .i_in(), .o_out(w2050135));
	wire w10136;
	torch #(1'b1) c10136 (.i_clk(tick), .i_in(), .o_out(w10136));
	wire w50136;
	torch #(1'b1) c50136 (.i_clk(tick), .i_in(), .o_out(w50136));
	wire w90136;
	torch #(1'b1) c90136 (.i_clk(tick), .i_in(), .o_out(w90136));
	wire w130136;
	torch #(1'b1) c130136 (.i_clk(tick), .i_in(), .o_out(w130136));
	wire w170136;
	torch #(1'b1) c170136 (.i_clk(tick), .i_in(), .o_out(w170136));
	wire w200136;
	repeater #(1, 1'b0, 0, 0) c200136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200136));
	wire w770136;
	repeater #(1, 1'b1, 0, 0) c770136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w770136));
	wire w1110136;
	repeater #(1, 1'b1, 0, 0) c1110136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1110136));
	wire w700137;
	repeater #(1, 1'b1, 0, 0) c700137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w700137));
	wire w830137;

	wire w860137;
	repeater #(1, 1'b1, 0, 0) c860137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w860137));
	wire w1040137;
	repeater #(1, 1'b1, 0, 0) c1040137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1040137));
	wire w1170137;

	wire w1200137;
	repeater #(1, 1'b1, 0, 0) c1200137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1200137));
	wire w750138;

	wire w1090138;

	wire w2000138;
	torch #(1'b0) c2000138 (.i_clk(tick), .i_in(), .o_out(w2000138));
	wire w2040138;
	torch #(1'b0) c2040138 (.i_clk(tick), .i_in(), .o_out(w2040138));
	wire w00139;
	torch #(1'b0) c00139 (.i_clk(tick), .i_in(), .o_out(w00139));
	wire w40139;
	torch #(1'b0) c40139 (.i_clk(tick), .i_in(), .o_out(w40139));
	wire w80139;
	torch #(1'b0) c80139 (.i_clk(tick), .i_in(), .o_out(w80139));
	wire w120139;
	torch #(1'b0) c120139 (.i_clk(tick), .i_in(), .o_out(w120139));
	wire w160139;
	torch #(1'b0) c160139 (.i_clk(tick), .i_in(), .o_out(w160139));
	wire w830139;

	wire w1170139;

	wire w700140;

	wire w800140;

	wire w850140;

	wire w860140;

	wire w1040140;

	wire w1140140;

	wire w1190140;

	wire w1200140;

	wire w620142;

	wire w690142;

	wire w780142;

	wire w960142;

	wire w1030142;

	wire w1120142;

	wire w840143;

	wire w850143;

	wire w1180143;

	wire w1190143;

	wire w780144;

	wire w1120144;

	wire w1390144;
	repeater #(2, 1'b1, 0, 0) c1390144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390144));
	wire w1410144;
	repeater #(1, 1'b1, 0, 0) c1410144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1410144));
	wire w1430144;
	repeater #(2, 1'b1, 0, 0) c1430144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1430144));
	wire w1450144;
	repeater #(1, 1'b0, 0, 0) c1450144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450144));
	wire w1470144;
	repeater #(2, 1'b1, 0, 0) c1470144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470144));
	wire w1490144;
	repeater #(1, 1'b1, 0, 0) c1490144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490144));
	wire w1510144;
	repeater #(2, 1'b1, 0, 0) c1510144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510144));
	wire w1530144;
	repeater #(1, 1'b1, 0, 0) c1530144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1530144));
	wire w1730144;
	repeater #(1, 1'b1, 0, 0) c1730144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1730144));
	wire w1750144;
	repeater #(2, 1'b1, 0, 0) c1750144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750144));
	wire w1770144;
	repeater #(1, 1'b1, 0, 0) c1770144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770144));
	wire w1790144;
	repeater #(2, 1'b1, 0, 0) c1790144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790144));
	wire w1810144;
	repeater #(1, 1'b0, 0, 0) c1810144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810144));
	wire w1830144;
	repeater #(2, 1'b1, 0, 0) c1830144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830144));
	wire w1850144;
	repeater #(1, 1'b1, 0, 0) c1850144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850144));
	wire w1870144;
	repeater #(2, 1'b1, 0, 0) c1870144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870144));
	wire w620146;

	wire w660146;

	wire w700146;

	wire w740146;

	wire w780146;

	wire w820146;

	wire w860146;

	wire w960146;

	wire w1000146;

	wire w1040146;

	wire w1080146;

	wire w1120146;

	wire w1160146;

	wire w1200146;

	wire w1480146;

	wire w1780146;

	wire w1400147;

	wire w1440147;

	wire w1470147;

	wire w1490147;

	wire w1520147;

	wire w1740147;

	wire w1770147;

	wire w1790147;

	wire w1820147;

	wire w1860147;

	wire w1390148;

	wire w1410148;

	wire w1430148;

	wire w1450148;

	wire w1480148;

	wire w1510148;

	wire w1530148;

	wire w1730148;

	wire w1750148;

	wire w1780148;

	wire w1810148;

	wire w1830148;

	wire w1850148;

	wire w1870148;

	wire w1440149;

	wire w1620149;
	repeater #(1, 1'b1, 0, 0) c1620149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620149));
	wire w1820149;

	wire w620150;

	wire w660150;

	wire w700150;

	wire w740150;

	wire w780150;

	wire w820150;

	wire w860150;

	wire w960150;

	wire w1000150;

	wire w1040150;

	wire w1080150;

	wire w1120150;

	wire w1160150;

	wire w1200150;

	wire w1400150;

	wire w1440150;

	wire w1450150;

	wire w1490150;

	wire w1510150;

	wire w1530150;

	wire w1730150;

	wire w1750150;

	wire w1770150;

	wire w1810150;

	wire w1820150;

	wire w1860150;

	wire w600152;
	repeater #(1, 1'b1, 0, 0) c600152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600152));
	wire w640152;
	repeater #(1, 1'b1, 0, 0) c640152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640152));
	wire w680152;
	repeater #(1, 1'b1, 0, 0) c680152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w680152));
	wire w720152;
	repeater #(1, 1'b1, 0, 0) c720152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w720152));
	wire w940152;
	repeater #(1, 1'b1, 0, 0) c940152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w940152));
	wire w980152;
	repeater #(1, 1'b1, 0, 0) c980152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w980152));
	wire w1020152;
	repeater #(1, 1'b1, 0, 0) c1020152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1020152));
	wire w1060152;
	repeater #(1, 1'b1, 0, 0) c1060152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060152));
	wire w1390152;

	wire w1450152;

	wire w1810152;

	wire w1870152;

	wire w780153;

	wire w820153;

	wire w860153;

	wire w1120153;

	wire w1160153;

	wire w1200153;

	wire w1350153;
	repeater #(1, 1'b1, 0, 0) c1350153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350153));
	wire w1400153;
	repeater #(1, 1'b1, 0, 0) c1400153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1400153));
	wire w1450153;
	repeater #(1, 1'b1, 0, 0) c1450153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450153));
	wire w1810153;
	repeater #(1, 1'b1, 0, 0) c1810153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810153));
	wire w1860153;
	repeater #(1, 1'b1, 0, 0) c1860153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860153));
	wire w1910153;
	repeater #(1, 1'b1, 0, 0) c1910153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910153));
	wire w2010153;
	torch #(1'b1) c2010153 (.i_clk(tick), .i_in(), .o_out(w2010153));
	wire w2050153;
	torch #(1'b1) c2050153 (.i_clk(tick), .i_in(), .o_out(w2050153));
	wire w10154;
	torch #(1'b1) c10154 (.i_clk(tick), .i_in(), .o_out(w10154));
	wire w50154;
	torch #(1'b1) c50154 (.i_clk(tick), .i_in(), .o_out(w50154));
	wire w90154;
	torch #(1'b1) c90154 (.i_clk(tick), .i_in(), .o_out(w90154));
	wire w130154;
	torch #(1'b1) c130154 (.i_clk(tick), .i_in(), .o_out(w130154));
	wire w170154;
	torch #(1'b1) c170154 (.i_clk(tick), .i_in(), .o_out(w170154));
	wire w2020154;
	repeater #(1, 1'b0, 0, 0) c2020154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020154));
	wire w2060154;
	repeater #(1, 1'b0, 0, 0) c2060154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060154));
	wire w20155;
	repeater #(1, 1'b0, 0, 0) c20155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20155));
	wire w60155;
	repeater #(1, 1'b0, 0, 0) c60155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60155));
	wire w100155;
	repeater #(1, 1'b0, 0, 0) c100155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100155));
	wire w140155;
	repeater #(1, 1'b0, 0, 0) c140155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140155));
	wire w180155;
	repeater #(1, 1'b0, 0, 0) c180155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180155));
	wire w780155;

	wire w1120155;

	wire w2000156;

	wire w2020156;
	repeater #(1, 1'b0, 0, 0) c2020156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020156));
	wire w2040156;

	wire w2060156;
	repeater #(1, 1'b0, 0, 0) c2060156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060156));
	wire w00157;

	wire w20157;
	repeater #(1, 1'b0, 0, 0) c20157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20157));
	wire w40157;

	wire w60157;
	repeater #(1, 1'b0, 0, 0) c60157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60157));
	wire w80157;

	wire w100157;
	repeater #(1, 1'b0, 0, 0) c100157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100157));
	wire w120157;

	wire w140157;
	repeater #(1, 1'b0, 0, 0) c140157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140157));
	wire w160157;

	wire w180157;
	repeater #(1, 1'b0, 0, 0) c180157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180157));
	wire w670157;
	repeater #(1, 1'b1, 0, 0) c670157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w670157));
	wire w700157;

	wire w830157;
	repeater #(1, 1'b0, 0, 0) c830157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w830157));
	wire w1010157;
	repeater #(1, 1'b1, 0, 0) c1010157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010157));
	wire w1040157;

	wire w1170157;
	repeater #(1, 1'b1, 0, 0) c1170157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1170157));
	wire w1340157;

	wire w1350157;
	repeater #(1, 1'b0, 0, 0) c1350157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350157));
	wire w1390157;

	wire w1400157;
	repeater #(1, 1'b0, 0, 0) c1400157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1400157));
	wire w1440157;

	wire w1450157;
	repeater #(1, 1'b1, 0, 0) c1450157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450157));
	wire w1810157;
	repeater #(1, 1'b1, 0, 0) c1810157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810157));
	wire w1820157;

	wire w1860157;
	repeater #(1, 1'b0, 0, 0) c1860157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860157));
	wire w1870157;

	wire w1910157;
	repeater #(1, 1'b1, 0, 0) c1910157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910157));
	wire w1920157;

	wire w780158;

	wire w1120158;

	wire w700159;

	wire w1040159;

	wire w670160;

	wire w680160;

	wire w730160;

	wire w810160;

	wire w830160;

	wire w1010160;

	wire w1020160;

	wire w1070160;

	wire w1150160;

	wire w1170160;

	wire w1350161;
	repeater #(2, 1'b0, 0, 0) c1350161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350161));
	wire w1400161;
	repeater #(2, 1'b0, 0, 0) c1400161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1400161));
	wire w1450161;
	repeater #(2, 1'b0, 0, 0) c1450161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1450161));
	wire w1810161;
	repeater #(2, 1'b1, 0, 0) c1810161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810161));
	wire w1860161;
	repeater #(2, 1'b0, 0, 0) c1860161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860161));
	wire w1910161;
	repeater #(2, 1'b0, 0, 0) c1910161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910161));
	wire w750162;

	wire w760162;

	wire w1090162;

	wire w1100162;

	wire w670164;

	wire w680164;

	wire w810164;

	wire w830164;

	wire w840164;

	wire w1010164;

	wire w1020164;

	wire w1150164;

	wire w1170164;

	wire w1180164;

	wire w780166;
	torch #(1'b1) c780166 (.i_clk(tick), .i_in(), .o_out(w780166));
	wire w790166;

	wire w1120166;
	torch #(1'b1) c1120166 (.i_clk(tick), .i_in(), .o_out(w1120166));
	wire w1130166;

	wire w1360166;
	repeater #(2, 1'b1, 0, 0) c1360166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1360166));
	wire w1630166;

	wire w1900166;
	repeater #(2, 1'b1, 0, 0) c1900166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1900166));
	wire w790167;

	wire w810167;

	wire w1130167;

	wire w1150167;

	wire w1340167;

	wire w1350167;

	wire w1410167;
	repeater #(1, 1'b0, 0, 0) c1410167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1410167));
	wire w1420167;
	repeater #(2, 1'b0, 0, 0) c1420167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420167));
	wire w1640167;

	wire w1840167;
	repeater #(2, 1'b1, 0, 0) c1840167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1840167));
	wire w1850167;
	repeater #(1, 1'b1, 0, 0) c1850167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850167));
	wire w1910167;

	wire w1920167;

	wire w1380168;
	repeater #(2, 1'b0, 0, 0) c1380168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380168));
	wire w1390168;
	repeater #(2, 1'b0, 0, 0) c1390168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390168));
	wire w1410168;

	wire w1550168;
	repeater #(1, 1'b0, 0, 0) c1550168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550168));
	wire w1560168;

	wire w1640168;
	repeater #(1, 1'b1, 0, 0) c1640168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640168));
	wire w1700168;

	wire w1710168;
	repeater #(1, 1'b0, 0, 0) c1710168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710168));
	wire w1850168;

	wire w1870168;
	repeater #(2, 1'b1, 0, 0) c1870168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870168));
	wire w1880168;
	repeater #(2, 1'b1, 0, 0) c1880168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1880168));
	wire w810169;

	wire w820169;

	wire w830169;

	wire w1150169;

	wire w1160169;

	wire w1170169;

	wire w1390169;

	wire w1410169;
	repeater #(1, 1'b1, 0, 0) c1410169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1410169));
	wire w1520169;

	wire w1530169;

	wire w1730169;

	wire w1740169;

	wire w1850169;
	repeater #(1, 1'b0, 0, 0) c1850169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850169));
	wire w1870169;

	wire w2010169;
	torch #(1'b1) c2010169 (.i_clk(tick), .i_in(), .o_out(w2010169));
	wire w2050169;
	torch #(1'b1) c2050169 (.i_clk(tick), .i_in(), .o_out(w2050169));
	wire w10170;
	torch #(1'b1) c10170 (.i_clk(tick), .i_in(), .o_out(w10170));
	wire w50170;
	torch #(1'b1) c50170 (.i_clk(tick), .i_in(), .o_out(w50170));
	wire w90170;
	torch #(1'b1) c90170 (.i_clk(tick), .i_in(), .o_out(w90170));
	wire w130170;
	torch #(1'b1) c130170 (.i_clk(tick), .i_in(), .o_out(w130170));
	wire w170170;
	torch #(1'b1) c170170 (.i_clk(tick), .i_in(), .o_out(w170170));
	wire w760170;

	wire w770170;

	wire w830170;

	wire w1100170;

	wire w1110170;

	wire w1170170;

	wire w1350170;

	wire w1390170;

	wire w1630170;

	wire w1640170;

	wire w1870170;

	wire w1910170;

	wire w2020170;
	repeater #(1, 1'b0, 0, 0) c2020170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020170));
	wire w2060170;
	repeater #(1, 1'b0, 0, 0) c2060170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060170));
	wire w20171;
	repeater #(1, 1'b0, 0, 0) c20171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20171));
	wire w60171;
	repeater #(1, 1'b0, 0, 0) c60171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60171));
	wire w100171;
	repeater #(1, 1'b0, 0, 0) c100171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100171));
	wire w140171;
	repeater #(1, 1'b0, 0, 0) c140171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140171));
	wire w180171;
	repeater #(1, 1'b0, 0, 0) c180171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180171));
	wire w1350171;

	wire w1370171;
	repeater #(1, 1'b0, 0, 0) c1370171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370171));
	wire w1420171;

	wire w1460171;

	wire w1520171;
	repeater #(1, 1'b0, 0, 0) c1520171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520171));
	wire w1600171;

	wire w1610171;
	repeater #(1, 1'b1, 0, 0) c1610171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610171));
	wire w1740171;
	repeater #(1, 1'b0, 0, 0) c1740171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1740171));
	wire w1800171;

	wire w1840171;

	wire w1890171;
	repeater #(1, 1'b1, 0, 0) c1890171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1890171));
	wire w1910171;

	wire w810172;
	repeater #(1, 1'b0, 0, 0) c810172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w810172));
	wire w830172;
	torch #(1'b0) c830172 (.i_clk(tick), .i_in(), .o_out(w830172));
	wire w890172;
	torch #(1'b1) c890172 (.i_clk(tick), .i_in(), .o_out(w890172));
	wire w1150172;
	repeater #(1, 1'b0, 0, 0) c1150172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1150172));
	wire w1170172;
	torch #(1'b0) c1170172 (.i_clk(tick), .i_in(), .o_out(w1170172));
	wire w1230172;
	torch #(1'b1) c1230172 (.i_clk(tick), .i_in(), .o_out(w1230172));
	wire w1420172;

	wire w1440172;
	repeater #(1, 1'b1, 0, 0) c1440172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1440172));
	wire w1450172;

	wire w1520172;

	wire w1690172;

	wire w1740172;

	wire w1810172;

	wire w1820172;
	repeater #(1, 1'b0, 0, 0) c1820172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820172));
	wire w1840172;

	wire w2000172;

	wire w2020172;
	repeater #(1, 1'b0, 0, 0) c2020172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020172));
	wire w2040172;

	wire w2060172;
	repeater #(1, 1'b0, 0, 0) c2060172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060172));
	wire w00173;

	wire w20173;
	repeater #(1, 1'b0, 0, 0) c20173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20173));
	wire w40173;

	wire w60173;
	repeater #(1, 1'b0, 0, 0) c60173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60173));
	wire w80173;

	wire w100173;
	repeater #(1, 1'b0, 0, 0) c100173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100173));
	wire w120173;

	wire w140173;
	repeater #(1, 1'b0, 0, 0) c140173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140173));
	wire w160173;

	wire w180173;
	repeater #(1, 1'b0, 0, 0) c180173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180173));
	wire w1380173;

	wire w1530173;

	wire w1570173;
	repeater #(1, 1'b0, 0, 0) c1570173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1570173));
	wire w1700173;
	repeater #(2, 1'b0, 0, 0) c1700173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1700173));
	wire w1730173;

	wire w1880173;

	wire w850174;
	repeater #(1, 1'b1, 0, 0) c850174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w850174));
	wire w1190174;
	repeater #(1, 1'b1, 0, 0) c1190174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190174));
	wire w1350174;

	wire w1360174;
	repeater #(1, 1'b0, 0, 0) c1360174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1360174));
	wire w1430174;
	repeater #(2, 1'b1, 0, 0) c1430174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1430174));
	wire w1560174;
	assign outputs[76] = ();
	wire w1830174;
	repeater #(2, 1'b0, 0, 0) c1830174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830174));
	wire w1900174;
	repeater #(1, 1'b0, 0, 0) c1900174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1900174));
	wire w1910174;

	wire w820176;
	torch #(1'b1) c820176 (.i_clk(tick), .i_in(), .o_out(w820176));
	wire w1160176;
	torch #(1'b1) c1160176 (.i_clk(tick), .i_in(), .o_out(w1160176));
	wire w900178;
	torch #(1'b1) c900178 (.i_clk(tick), .i_in(), .o_out(w900178));
	wire w1240178;
	torch #(1'b1) c1240178 (.i_clk(tick), .i_in(), .o_out(w1240178));
	wire w8110;
	repeater #(2, 1'b0, 0, 0) c8110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8110));
	wire w11510;
	repeater #(2, 1'b0, 0, 0) c11510 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11510));
	wire w9111;
	repeater #(2, 1'b0, 0, 0) c9111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9111));
	wire w12511;
	repeater #(2, 1'b0, 0, 0) c12511 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12511));
	wire w6914;
	torch #(1'b0) c6914 (.i_clk(tick), .i_in(), .o_out(w6914));
	wire w7014;
	torch #(1'b0) c7014 (.i_clk(tick), .i_in(), .o_out(w7014));
	wire w7714;
	torch #(1'b0) c7714 (.i_clk(tick), .i_in(), .o_out(w7714));
	wire w7814;
	torch #(1'b0) c7814 (.i_clk(tick), .i_in(), .o_out(w7814));
	wire w8514;
	torch #(1'b0) c8514 (.i_clk(tick), .i_in(), .o_out(w8514));
	wire w8614;
	torch #(1'b0) c8614 (.i_clk(tick), .i_in(), .o_out(w8614));
	wire w10314;
	torch #(1'b0) c10314 (.i_clk(tick), .i_in(), .o_out(w10314));
	wire w10414;
	torch #(1'b0) c10414 (.i_clk(tick), .i_in(), .o_out(w10414));
	wire w11114;
	torch #(1'b0) c11114 (.i_clk(tick), .i_in(), .o_out(w11114));
	wire w11214;
	torch #(1'b0) c11214 (.i_clk(tick), .i_in(), .o_out(w11214));
	wire w11914;
	torch #(1'b0) c11914 (.i_clk(tick), .i_in(), .o_out(w11914));
	wire w12014;
	torch #(1'b0) c12014 (.i_clk(tick), .i_in(), .o_out(w12014));
	wire w6616;
	torch #(1'b1) c6616 (.i_clk(tick), .i_in(), .o_out(w6616));
	wire w6816;
	torch #(1'b1) c6816 (.i_clk(tick), .i_in(), .o_out(w6816));
	wire w7316;
	torch #(1'b1) c7316 (.i_clk(tick), .i_in(), .o_out(w7316));
	wire w7616;
	torch #(1'b1) c7616 (.i_clk(tick), .i_in(), .o_out(w7616));
	wire w8116;
	torch #(1'b1) c8116 (.i_clk(tick), .i_in(), .o_out(w8116));
	wire w8416;
	torch #(1'b1) c8416 (.i_clk(tick), .i_in(), .o_out(w8416));
	wire w8916;
	torch #(1'b1) c8916 (.i_clk(tick), .i_in(), .o_out(w8916));
	wire w10016;
	torch #(1'b1) c10016 (.i_clk(tick), .i_in(), .o_out(w10016));
	wire w10216;
	torch #(1'b1) c10216 (.i_clk(tick), .i_in(), .o_out(w10216));
	wire w10716;
	torch #(1'b1) c10716 (.i_clk(tick), .i_in(), .o_out(w10716));
	wire w11016;
	torch #(1'b1) c11016 (.i_clk(tick), .i_in(), .o_out(w11016));
	wire w11516;
	torch #(1'b1) c11516 (.i_clk(tick), .i_in(), .o_out(w11516));
	wire w11816;
	torch #(1'b1) c11816 (.i_clk(tick), .i_in(), .o_out(w11816));
	wire w12316;
	torch #(1'b1) c12316 (.i_clk(tick), .i_in(), .o_out(w12316));
	wire w20116;
	torch #(1'b1) c20116 (.i_clk(tick), .i_in(), .o_out(w20116));
	wire w20516;
	torch #(1'b1) c20516 (.i_clk(tick), .i_in(), .o_out(w20516));
	wire w117;
	torch #(1'b1) c117 (.i_clk(tick), .i_in(), .o_out(w117));
	wire w517;
	torch #(1'b1) c517 (.i_clk(tick), .i_in(), .o_out(w517));
	wire w917;
	torch #(1'b1) c917 (.i_clk(tick), .i_in(), .o_out(w917));
	wire w1317;
	torch #(1'b1) c1317 (.i_clk(tick), .i_in(), .o_out(w1317));
	wire w1717;
	torch #(1'b1) c1717 (.i_clk(tick), .i_in(), .o_out(w1717));
	wire w20217;
	repeater #(1, 1'b0, 0, 0) c20217 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20217));
	wire w20617;
	repeater #(1, 1'b0, 0, 0) c20617 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20617));
	wire w218;
	repeater #(1, 1'b0, 0, 0) c218 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w218));
	wire w618;
	repeater #(1, 1'b0, 0, 0) c618 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w618));
	wire w1018;
	repeater #(1, 1'b0, 0, 0) c1018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1018));
	wire w1418;
	repeater #(1, 1'b0, 0, 0) c1418 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1418));
	wire w1818;
	repeater #(1, 1'b0, 0, 0) c1818 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1818));
	wire w7718;
	repeater #(2, 1'b0, 0, 0) c7718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7718));
	wire w11118;
	repeater #(2, 1'b0, 0, 0) c11118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11118));
	wire w7719;
	repeater #(1, 1'b0, 0, 0) c7719 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7719));
	wire w11119;
	repeater #(1, 1'b0, 0, 0) c11119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11119));
	wire w20019;

	wire w20219;
	repeater #(1, 1'b0, 0, 0) c20219 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20219));
	wire w20419;

	wire w20619;
	repeater #(1, 1'b0, 0, 0) c20619 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20619));
	wire w0110;

	wire w2110;
	repeater #(1, 1'b0, 0, 0) c2110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2110));
	wire w4110;

	wire w6110;
	repeater #(1, 1'b0, 0, 0) c6110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6110));
	wire w8110;

	wire w10110;
	repeater #(1, 1'b0, 0, 0) c10110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10110));
	wire w12110;

	wire w14110;
	repeater #(1, 1'b0, 0, 0) c14110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14110));
	wire w16110;

	wire w18110;
	repeater #(1, 1'b0, 0, 0) c18110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18110));
	wire w95110;
	repeater #(1, 1'b0, 0, 0) c95110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95110));
	wire w111110;
	repeater #(1, 1'b0, 0, 0) c111110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111110));
	wire w162117;

	wire w163117;
	repeater #(1, 1'b0, 0, 0) c163117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163117));
	wire w164118;
	repeater #(1, 1'b0, 0, 0) c164118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164118));
	wire w167118;
	repeater #(2, 1'b0, 0, 0) c167118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167118));
	wire w159119;
	repeater #(1, 1'b0, 0, 0) c159119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159119));
	wire w172119;
	repeater #(2, 1'b0, 0, 0) c172119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172119));
	wire w158120;
	assign outputs[77] = ();
	wire w161120;

	wire w170120;

	wire w161121;

	wire w170121;

	wire w159122;
	repeater #(1, 1'b0, 0, 0) c159122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159122));
	wire w172122;
	repeater #(1, 1'b0, 0, 0) c172122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172122));
	wire w201122;
	torch #(1'b1) c201122 (.i_clk(tick), .i_in(), .o_out(w201122));
	wire w205122;
	torch #(1'b1) c205122 (.i_clk(tick), .i_in(), .o_out(w205122));
	wire w1123;
	torch #(1'b1) c1123 (.i_clk(tick), .i_in(), .o_out(w1123));
	wire w5123;
	torch #(1'b1) c5123 (.i_clk(tick), .i_in(), .o_out(w5123));
	wire w9123;
	torch #(1'b1) c9123 (.i_clk(tick), .i_in(), .o_out(w9123));
	wire w13123;
	torch #(1'b1) c13123 (.i_clk(tick), .i_in(), .o_out(w13123));
	wire w17123;
	torch #(1'b1) c17123 (.i_clk(tick), .i_in(), .o_out(w17123));
	wire w202123;
	repeater #(1, 1'b0, 0, 0) c202123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202123));
	wire w206123;
	repeater #(1, 1'b0, 0, 0) c206123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206123));
	wire w2124;
	repeater #(1, 1'b0, 0, 0) c2124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2124));
	wire w6124;
	repeater #(1, 1'b0, 0, 0) c6124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6124));
	wire w10124;
	repeater #(1, 1'b0, 0, 0) c10124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10124));
	wire w14124;
	repeater #(1, 1'b0, 0, 0) c14124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14124));
	wire w18124;
	repeater #(1, 1'b0, 0, 0) c18124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18124));
	wire w200125;

	wire w202125;
	repeater #(1, 1'b0, 0, 0) c202125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202125));
	wire w204125;

	wire w206125;
	repeater #(1, 1'b0, 0, 0) c206125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206125));
	wire w0126;

	wire w2126;
	repeater #(1, 1'b0, 0, 0) c2126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2126));
	wire w4126;

	wire w6126;
	repeater #(1, 1'b0, 0, 0) c6126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6126));
	wire w8126;

	wire w10126;
	repeater #(1, 1'b0, 0, 0) c10126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10126));
	wire w12126;

	wire w14126;
	repeater #(1, 1'b0, 0, 0) c14126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14126));
	wire w16126;

	wire w18126;
	repeater #(1, 1'b0, 0, 0) c18126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18126));
	wire w201138;
	torch #(1'b1) c201138 (.i_clk(tick), .i_in(), .o_out(w201138));
	wire w205138;
	torch #(1'b1) c205138 (.i_clk(tick), .i_in(), .o_out(w205138));
	wire w1139;
	torch #(1'b1) c1139 (.i_clk(tick), .i_in(), .o_out(w1139));
	wire w5139;
	torch #(1'b1) c5139 (.i_clk(tick), .i_in(), .o_out(w5139));
	wire w9139;
	torch #(1'b1) c9139 (.i_clk(tick), .i_in(), .o_out(w9139));
	wire w13139;
	torch #(1'b1) c13139 (.i_clk(tick), .i_in(), .o_out(w13139));
	wire w17139;
	torch #(1'b1) c17139 (.i_clk(tick), .i_in(), .o_out(w17139));
	wire w202139;
	repeater #(1, 1'b0, 0, 0) c202139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202139));
	wire w206139;
	repeater #(1, 1'b0, 0, 0) c206139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206139));
	wire w2140;
	repeater #(1, 1'b0, 0, 0) c2140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2140));
	wire w6140;
	repeater #(1, 1'b0, 0, 0) c6140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6140));
	wire w10140;
	repeater #(1, 1'b0, 0, 0) c10140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10140));
	wire w14140;
	repeater #(1, 1'b0, 0, 0) c14140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14140));
	wire w18140;
	repeater #(1, 1'b0, 0, 0) c18140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18140));
	wire w200141;

	wire w202141;
	repeater #(1, 1'b0, 0, 0) c202141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202141));
	wire w204141;

	wire w206141;
	repeater #(1, 1'b0, 0, 0) c206141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206141));
	wire w0142;

	wire w2142;
	repeater #(1, 1'b0, 0, 0) c2142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2142));
	wire w4142;

	wire w6142;
	repeater #(1, 1'b0, 0, 0) c6142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6142));
	wire w8142;

	wire w10142;
	repeater #(1, 1'b0, 0, 0) c10142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10142));
	wire w12142;

	wire w14142;
	repeater #(1, 1'b0, 0, 0) c14142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14142));
	wire w16142;

	wire w18142;
	repeater #(1, 1'b0, 0, 0) c18142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18142));
	wire w201147;
	torch #(1'b1) c201147 (.i_clk(tick), .i_in(), .o_out(w201147));
	wire w205147;
	torch #(1'b1) c205147 (.i_clk(tick), .i_in(), .o_out(w205147));
	wire w1148;
	torch #(1'b1) c1148 (.i_clk(tick), .i_in(), .o_out(w1148));
	wire w5148;
	torch #(1'b1) c5148 (.i_clk(tick), .i_in(), .o_out(w5148));
	wire w9148;
	torch #(1'b1) c9148 (.i_clk(tick), .i_in(), .o_out(w9148));
	wire w13148;
	torch #(1'b1) c13148 (.i_clk(tick), .i_in(), .o_out(w13148));
	wire w17148;
	torch #(1'b1) c17148 (.i_clk(tick), .i_in(), .o_out(w17148));
	wire w201156;
	repeater #(1, 1'b0, 0, 0) c201156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201156));
	wire w205156;
	repeater #(1, 1'b0, 0, 0) c205156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205156));
	wire w1157;
	repeater #(1, 1'b0, 0, 0) c1157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1157));
	wire w5157;
	repeater #(1, 1'b0, 0, 0) c5157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5157));
	wire w9157;
	repeater #(1, 1'b0, 0, 0) c9157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9157));
	wire w13157;
	repeater #(1, 1'b0, 0, 0) c13157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13157));
	wire w17157;
	repeater #(1, 1'b0, 0, 0) c17157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17157));
	wire w202159;
	repeater #(1, 1'b0, 0, 0) c202159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202159));
	wire w206159;
	repeater #(1, 1'b0, 0, 0) c206159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206159));
	wire w2160;
	repeater #(1, 1'b0, 0, 0) c2160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2160));
	wire w6160;
	repeater #(1, 1'b0, 0, 0) c6160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6160));
	wire w10160;
	repeater #(1, 1'b0, 0, 0) c10160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10160));
	wire w14160;
	repeater #(1, 1'b0, 0, 0) c14160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14160));
	wire w18160;
	repeater #(1, 1'b0, 0, 0) c18160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18160));
	wire w201160;
	repeater #(1, 1'b1, 0, 0) c201160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201160));
	wire w205160;
	repeater #(1, 1'b1, 0, 0) c205160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205160));
	wire w1161;
	repeater #(1, 1'b1, 0, 0) c1161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161));
	wire w5161;
	repeater #(1, 1'b0, 0, 0) c5161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5161));
	wire w9161;
	repeater #(1, 1'b1, 0, 0) c9161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9161));
	wire w13161;
	repeater #(1, 1'b1, 0, 0) c13161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13161));
	wire w17161;
	repeater #(1, 1'b1, 0, 0) c17161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17161));
	wire w201194;
	torch #(1'b1) c201194 (.i_clk(tick), .i_in(), .o_out(w201194));
	wire w205194;
	torch #(1'b1) c205194 (.i_clk(tick), .i_in(), .o_out(w205194));
	wire w1195;
	torch #(1'b1) c1195 (.i_clk(tick), .i_in(), .o_out(w1195));
	wire w5195;
	torch #(1'b1) c5195 (.i_clk(tick), .i_in(), .o_out(w5195));
	wire w9195;
	torch #(1'b1) c9195 (.i_clk(tick), .i_in(), .o_out(w9195));
	wire w13195;
	torch #(1'b1) c13195 (.i_clk(tick), .i_in(), .o_out(w13195));
	wire w17195;
	torch #(1'b1) c17195 (.i_clk(tick), .i_in(), .o_out(w17195));
	wire w109199;

	wire w143199;

	wire w177199;

	wire w31100;

	wire w1081100;
	repeater #(1, 1'b1, 0, 0) c1081100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081100));
	wire w1421100;
	repeater #(1, 1'b1, 0, 0) c1421100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1421100));
	wire w1761100;
	repeater #(1, 1'b1, 0, 0) c1761100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1761100));
	wire w21101;
	repeater #(1, 1'b1, 0, 0) c21101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21101));
	wire w1071101;

	wire w1411101;

	wire w1751101;

	wire w11102;

	wire w1061102;
	repeater #(1, 1'b0, 0, 0) c1061102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061102));
	wire w1401102;
	repeater #(1, 1'b0, 0, 0) c1401102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401102));
	wire w1741102;
	repeater #(1, 1'b1, 0, 0) c1741102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741102));
	wire w01103;
	repeater #(1, 1'b1, 0, 0) c01103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w01103));
	wire w1051103;

	wire w1391103;

	wire w1731103;

	wire w2071103;

	wire w1041104;
	repeater #(1, 1'b1, 0, 0) c1041104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1041104));
	wire w1381104;
	repeater #(1, 1'b1, 0, 0) c1381104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1381104));
	wire w1721104;
	repeater #(1, 1'b1, 0, 0) c1721104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1721104));
	wire w2061104;
	repeater #(1, 1'b1, 0, 0) c2061104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2061104));
	wire w1031105;

	wire w1371105;

	wire w1711105;

	wire w2051105;

	wire w1021106;
	repeater #(1, 1'b1, 0, 0) c1021106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1021106));
	wire w1361106;
	repeater #(1, 1'b1, 0, 0) c1361106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361106));
	wire w1701106;
	repeater #(1, 1'b1, 0, 0) c1701106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701106));
	wire w2041106;
	repeater #(1, 1'b1, 0, 0) c2041106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2041106));
	wire w1011107;

	wire w1351107;

	wire w1691107;

	wire w2031107;

	wire w1001108;
	repeater #(1, 1'b1, 0, 0) c1001108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1001108));
	wire w1341108;
	repeater #(1, 1'b1, 0, 0) c1341108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1341108));
	wire w1681108;
	repeater #(1, 1'b1, 0, 0) c1681108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1681108));
	wire w2021108;
	repeater #(1, 1'b1, 0, 0) c2021108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021108));
	wire w991109;

	wire w1331109;

	wire w1671109;

	wire w2011109;

	wire w981110;
	repeater #(1, 1'b1, 0, 0) c981110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981110));
	wire w1321110;
	repeater #(1, 1'b1, 0, 0) c1321110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321110));
	wire w1661110;
	repeater #(1, 1'b1, 0, 0) c1661110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661110));
	wire w2001110;
	repeater #(1, 1'b1, 0, 0) c2001110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2001110));
	wire w971111;

	wire w1311111;

	wire w1651111;

	wire w1991111;

	wire w961112;
	repeater #(1, 1'b1, 0, 0) c961112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w961112));
	wire w1301112;
	repeater #(1, 1'b1, 0, 0) c1301112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1301112));
	wire w1641112;
	repeater #(1, 1'b1, 0, 0) c1641112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1641112));
	wire w1981112;
	repeater #(1, 1'b1, 0, 0) c1981112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1981112));
	wire w951113;

	wire w1291113;

	wire w1631113;

	wire w1971113;

	wire w941114;
	repeater #(1, 1'b1, 0, 0) c941114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941114));
	wire w1281114;
	repeater #(1, 1'b1, 0, 0) c1281114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281114));
	wire w1621114;
	repeater #(1, 1'b1, 0, 0) c1621114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621114));
	wire w1961114;
	repeater #(1, 1'b1, 0, 0) c1961114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1961114));
	wire w931115;

	wire w1271115;

	wire w1611115;

	wire w1951115;

	wire w921116;
	repeater #(1, 1'b1, 0, 0) c921116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w921116));
	wire w1261116;
	repeater #(1, 1'b1, 0, 0) c1261116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1261116));
	wire w1601116;
	repeater #(1, 1'b1, 0, 0) c1601116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1601116));
	wire w1941116;
	repeater #(1, 1'b1, 0, 0) c1941116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941116));
	wire w911117;

	wire w1251117;

	wire w1591117;

	wire w1931117;

	wire w901118;
	repeater #(1, 1'b1, 0, 0) c901118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901118));
	wire w1241118;
	repeater #(1, 1'b1, 0, 0) c1241118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241118));
	wire w1581118;
	repeater #(1, 1'b1, 0, 0) c1581118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581118));
	wire w1921118;
	repeater #(1, 1'b1, 0, 0) c1921118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1921118));
	wire w891119;

	wire w1231119;

	wire w1571119;

	wire w1911119;

	wire w881120;
	repeater #(1, 1'b1, 0, 0) c881120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w881120));
	wire w1221120;
	repeater #(1, 1'b1, 0, 0) c1221120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1221120));
	wire w1561120;
	repeater #(1, 1'b1, 0, 0) c1561120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1561120));
	wire w1901120;
	repeater #(1, 1'b1, 0, 0) c1901120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901120));
	wire w871121;

	wire w1211121;

	wire w1551121;

	wire w1891121;

	wire w861122;
	repeater #(1, 1'b1, 0, 0) c861122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861122));
	wire w1201122;
	repeater #(1, 1'b1, 0, 0) c1201122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201122));
	wire w1541122;
	repeater #(1, 1'b1, 0, 0) c1541122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541122));
	wire w1881122;
	repeater #(1, 1'b1, 0, 0) c1881122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1881122));
	wire w851123;

	wire w1191123;

	wire w1531123;

	wire w1871123;

	wire w841124;
	repeater #(1, 1'b1, 0, 0) c841124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w841124));
	wire w1181124;
	repeater #(1, 1'b1, 0, 0) c1181124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1181124));
	wire w1521124;
	repeater #(1, 1'b1, 0, 0) c1521124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1521124));
	wire w1861124;
	repeater #(1, 1'b1, 0, 0) c1861124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861124));
	wire w831125;

	wire w1171125;

	wire w1511125;

	wire w1851125;

	wire w821126;
	repeater #(1, 1'b1, 0, 0) c821126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821126));
	wire w1161126;
	repeater #(1, 1'b1, 0, 0) c1161126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161126));
	wire w1501126;
	repeater #(1, 1'b1, 0, 0) c1501126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1501126));
	wire w1841126;
	repeater #(1, 1'b1, 0, 0) c1841126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1841126));
	wire w1331130;
	torch #(1'b0) c1331130 (.i_clk(tick), .i_in(), .o_out(w1331130));
	wire w1371130;
	torch #(1'b0) c1371130 (.i_clk(tick), .i_in(), .o_out(w1371130));
	wire w1411130;
	torch #(1'b0) c1411130 (.i_clk(tick), .i_in(), .o_out(w1411130));
	wire w1451130;
	torch #(1'b1) c1451130 (.i_clk(tick), .i_in(), .o_out(w1451130));
	wire w1491130;
	torch #(1'b0) c1491130 (.i_clk(tick), .i_in(), .o_out(w1491130));
	wire w1531130;
	torch #(1'b0) c1531130 (.i_clk(tick), .i_in(), .o_out(w1531130));
	wire w1571130;
	torch #(1'b0) c1571130 (.i_clk(tick), .i_in(), .o_out(w1571130));
	wire w1691130;
	torch #(1'b0) c1691130 (.i_clk(tick), .i_in(), .o_out(w1691130));
	wire w1731130;
	torch #(1'b0) c1731130 (.i_clk(tick), .i_in(), .o_out(w1731130));
	wire w1771130;
	torch #(1'b0) c1771130 (.i_clk(tick), .i_in(), .o_out(w1771130));
	wire w1811130;
	torch #(1'b1) c1811130 (.i_clk(tick), .i_in(), .o_out(w1811130));
	wire w1851130;
	torch #(1'b0) c1851130 (.i_clk(tick), .i_in(), .o_out(w1851130));
	wire w1891130;
	torch #(1'b0) c1891130 (.i_clk(tick), .i_in(), .o_out(w1891130));
	wire w1931130;
	torch #(1'b0) c1931130 (.i_clk(tick), .i_in(), .o_out(w1931130));
	wire w801131;
	repeater #(2, 1'b1, 0, 0) c801131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w801131));
	wire w1141131;
	repeater #(2, 1'b1, 0, 0) c1141131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1141131));
	wire w2001132;
	repeater #(1, 1'b1, 0, 0) c2001132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2001132));
	wire w2041132;
	repeater #(1, 1'b1, 0, 0) c2041132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2041132));
	wire w01133;
	repeater #(1, 1'b1, 0, 0) c01133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w01133));
	wire w41133;
	repeater #(1, 1'b1, 0, 0) c41133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41133));
	wire w81133;
	repeater #(1, 1'b1, 0, 0) c81133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81133));
	wire w121133;
	repeater #(1, 1'b1, 0, 0) c121133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121133));
	wire w161133;
	repeater #(1, 1'b1, 0, 0) c161133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161133));
	wire w661133;
	repeater #(1, 1'b1, 0, 0) c661133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w661133));
	wire w721133;
	torch #(1'b1) c721133 (.i_clk(tick), .i_in(), .o_out(w721133));
	wire w821133;
	repeater #(1, 1'b1, 0, 0) c821133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821133));
	wire w1001133;
	repeater #(1, 1'b1, 0, 0) c1001133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1001133));
	wire w1061133;
	torch #(1'b1) c1061133 (.i_clk(tick), .i_in(), .o_out(w1061133));
	wire w1161133;
	repeater #(1, 1'b1, 0, 0) c1161133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161133));
	wire w2001133;
	repeater #(1, 1'b1, 0, 0) c2001133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2001133));
	wire w2021133;
	repeater #(1, 1'b0, 0, 0) c2021133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021133));
	wire w2041133;
	repeater #(1, 1'b1, 0, 0) c2041133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2041133));
	wire w2061133;
	repeater #(1, 1'b0, 0, 0) c2061133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2061133));
	wire w01134;
	repeater #(1, 1'b1, 0, 0) c01134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w01134));
	wire w21134;
	repeater #(1, 1'b0, 0, 0) c21134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21134));
	wire w41134;
	repeater #(1, 1'b1, 0, 0) c41134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41134));
	wire w61134;
	repeater #(1, 1'b0, 0, 0) c61134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61134));
	wire w81134;
	repeater #(1, 1'b1, 0, 0) c81134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81134));
	wire w101134;
	repeater #(1, 1'b0, 0, 0) c101134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101134));
	wire w121134;
	repeater #(1, 1'b1, 0, 0) c121134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121134));
	wire w141134;
	repeater #(1, 1'b0, 0, 0) c141134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141134));
	wire w161134;
	repeater #(1, 1'b1, 0, 0) c161134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161134));
	wire w181134;
	repeater #(1, 1'b0, 0, 0) c181134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w181134));
	wire w2011134;
	torch #(1'b0) c2011134 (.i_clk(tick), .i_in(), .o_out(w2011134));
	wire w2051134;
	torch #(1'b0) c2051134 (.i_clk(tick), .i_in(), .o_out(w2051134));
	wire w11135;
	torch #(1'b0) c11135 (.i_clk(tick), .i_in(), .o_out(w11135));
	wire w51135;
	torch #(1'b0) c51135 (.i_clk(tick), .i_in(), .o_out(w51135));
	wire w91135;
	torch #(1'b0) c91135 (.i_clk(tick), .i_in(), .o_out(w91135));
	wire w131135;
	torch #(1'b0) c131135 (.i_clk(tick), .i_in(), .o_out(w131135));
	wire w171135;
	torch #(1'b0) c171135 (.i_clk(tick), .i_in(), .o_out(w171135));
	wire w5001;
	repeater #(1, 1'b1, 0, 0) c5001 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5001));
	wire w6301;

	wire w6601;
	repeater #(1, 1'b1, 0, 0) c6601 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6601));
	wire w8401;
	repeater #(1, 1'b1, 0, 0) c8401 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8401));
	wire w9701;

	wire w10001;
	repeater #(1, 1'b1, 0, 0) c10001 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10001));
	wire w11701;
	repeater #(1, 1'b1, 0, 0) c11701 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11701));
	wire w12101;
	repeater #(1, 1'b1, 0, 0) c12101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12101));
	wire w12501;
	repeater #(1, 1'b1, 0, 0) c12501 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12501));
	wire w12901;
	repeater #(1, 1'b0, 0, 0) c12901 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12901));
	wire w13301;
	repeater #(1, 1'b1, 0, 0) c13301 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13301));
	wire w13701;
	repeater #(1, 1'b1, 0, 0) c13701 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13701));
	wire w14101;
	repeater #(1, 1'b1, 0, 0) c14101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14101));
	wire w15301;
	repeater #(1, 1'b1, 0, 0) c15301 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15301));
	wire w15701;
	repeater #(1, 1'b1, 0, 0) c15701 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15701));
	wire w16101;
	repeater #(1, 1'b1, 0, 0) c16101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16101));
	wire w16501;
	repeater #(1, 1'b0, 0, 0) c16501 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16501));
	wire w16901;
	repeater #(1, 1'b1, 0, 0) c16901 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16901));
	wire w17301;
	repeater #(1, 1'b1, 0, 0) c17301 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17301));
	wire w17701;
	repeater #(1, 1'b1, 0, 0) c17701 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17701));
	wire w5502;

	wire w8902;

	wire w6303;

	wire w9703;

	wire w5004;

	wire w6004;

	wire w6504;

	wire w6604;

	wire w8404;

	wire w9404;

	wire w9904;

	wire w10004;

	wire w5806;

	wire w9206;

	wire w4907;

	wire w6407;

	wire w6507;

	wire w8307;

	wire w9807;

	wire w9907;

	wire w5008;

	wire w5408;

	wire w5808;

	wire w8408;

	wire w8808;

	wire w9208;

	wire w18608;

	wire w19008;

	wire w19408;

	wire w19808;

	wire w20208;

	wire w20608;

	wire w209;

	wire w74011;

	wire w108011;

	wire w47012;

	wire w48012;

	wire w51012;

	wire w52012;

	wire w55012;

	wire w56012;

	wire w59012;

	wire w60012;

	wire w63012;

	wire w64012;

	wire w67012;

	wire w68012;

	wire w71012;

	wire w72012;

	wire w81012;

	wire w82012;

	wire w85012;

	wire w86012;

	wire w89012;

	wire w90012;

	wire w93012;

	wire w94012;

	wire w97012;

	wire w98012;

	wire w101012;

	wire w102012;

	wire w105012;

	wire w106012;

	wire w145012;

	wire w45013;

	wire w79013;

	wire w60016;
	repeater #(1, 1'b1, 0, 0) c60016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60016));
	wire w64016;
	repeater #(1, 1'b1, 0, 0) c64016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64016));
	wire w68016;
	repeater #(1, 1'b1, 0, 0) c68016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68016));
	wire w94016;
	repeater #(1, 1'b1, 0, 0) c94016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94016));
	wire w98016;
	repeater #(1, 1'b1, 0, 0) c98016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98016));
	wire w102016;
	repeater #(1, 1'b1, 0, 0) c102016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102016));
	wire w66019;

	wire w70019;

	wire w100019;

	wire w104019;

	wire w186019;
	torch #(1'b0) c186019 (.i_clk(tick), .i_in(), .o_out(w186019));
	wire w190019;
	torch #(1'b0) c190019 (.i_clk(tick), .i_in(), .o_out(w190019));
	wire w194019;
	torch #(1'b0) c194019 (.i_clk(tick), .i_in(), .o_out(w194019));
	wire w198019;
	torch #(1'b0) c198019 (.i_clk(tick), .i_in(), .o_out(w198019));
	wire w202019;
	torch #(1'b0) c202019 (.i_clk(tick), .i_in(), .o_out(w202019));
	wire w206019;
	torch #(1'b0) c206019 (.i_clk(tick), .i_in(), .o_out(w206019));
	wire w2020;
	torch #(1'b0) c2020 (.i_clk(tick), .i_in(), .o_out(w2020));
	wire w118020;
	repeater #(2, 1'b0, 0, 0) c118020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118020));
	wire w123020;
	repeater #(2, 1'b0, 0, 0) c123020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123020));
	wire w128020;
	repeater #(2, 1'b1, 0, 0) c128020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128020));
	wire w166020;
	repeater #(2, 1'b1, 0, 0) c166020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166020));
	wire w171020;
	repeater #(2, 1'b0, 0, 0) c171020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171020));
	wire w176020;
	repeater #(2, 1'b1, 0, 0) c176020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176020));
	wire w55021;
	repeater #(1, 1'b1, 0, 0) c55021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55021));
	wire w89021;
	repeater #(1, 1'b1, 0, 0) c89021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89021));
	wire w66022;

	wire w100022;

	wire w55024;

	wire w56024;

	wire w69024;

	wire w89024;

	wire w90024;

	wire w103024;

	wire w186024;

	wire w190024;

	wire w194024;

	wire w198024;

	wire w202024;

	wire w206024;

	wire w2025;

	wire w55028;

	wire w56028;

	wire w69028;

	wire w89028;

	wire w90028;

	wire w103028;

	wire w145029;
	assign outputs[78] = ();
	wire w66030;
	torch #(1'b1) c66030 (.i_clk(tick), .i_in(), .o_out(w66030));
	wire w67030;

	wire w100030;
	torch #(1'b1) c100030 (.i_clk(tick), .i_in(), .o_out(w100030));
	wire w101030;

	wire w67031;

	wire w69031;

	wire w101031;

	wire w103031;

	wire w117031;
	repeater #(1, 1'b0, 0, 0) c117031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117031));
	wire w149031;

	wire w177031;
	repeater #(1, 1'b1, 0, 0) c177031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177031));
	wire w121032;
	repeater #(1, 1'b0, 0, 0) c121032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121032));
	wire w146032;

	wire w173032;
	repeater #(1, 1'b1, 0, 0) c173032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173032));
	wire w69033;

	wire w70033;

	wire w71033;

	wire w103033;

	wire w104033;

	wire w105033;

	wire w127033;

	wire w131033;
	repeater #(1, 1'b1, 0, 0) c131033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131033));
	wire w145033;

	wire w147033;
	repeater #(2, 1'b1, 0, 0) c147033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147033));
	wire w150033;
	repeater #(2, 1'b1, 0, 0) c150033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150033));
	wire w163033;
	repeater #(1, 1'b1, 0, 0) c163033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163033));
	wire w167033;

	wire w64034;

	wire w65034;

	wire w71034;

	wire w98034;

	wire w99034;

	wire w105034;

	wire w128034;

	wire w134034;
	repeater #(2, 1'b0, 0, 0) c134034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134034));
	wire w137034;
	repeater #(2, 1'b0, 0, 0) c137034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137034));
	wire w139034;

	wire w155034;

	wire w157034;
	repeater #(2, 1'b0, 0, 0) c157034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157034));
	wire w160034;
	repeater #(2, 1'b0, 0, 0) c160034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160034));
	wire w166034;

	wire w127035;
	repeater #(2, 1'b0, 0, 0) c127035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127035));
	wire w138035;

	wire w156035;

	wire w167035;
	repeater #(2, 1'b1, 0, 0) c167035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167035));
	wire w186035;
	torch #(1'b0) c186035 (.i_clk(tick), .i_in(), .o_out(w186035));
	wire w190035;
	torch #(1'b0) c190035 (.i_clk(tick), .i_in(), .o_out(w190035));
	wire w194035;
	torch #(1'b0) c194035 (.i_clk(tick), .i_in(), .o_out(w194035));
	wire w198035;
	torch #(1'b0) c198035 (.i_clk(tick), .i_in(), .o_out(w198035));
	wire w202035;
	torch #(1'b0) c202035 (.i_clk(tick), .i_in(), .o_out(w202035));
	wire w206035;
	torch #(1'b0) c206035 (.i_clk(tick), .i_in(), .o_out(w206035));
	wire w2036;
	torch #(1'b0) c2036 (.i_clk(tick), .i_in(), .o_out(w2036));
	wire w69036;
	repeater #(1, 1'b0, 0, 0) c69036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69036));
	wire w71036;
	torch #(1'b0) c71036 (.i_clk(tick), .i_in(), .o_out(w71036));
	wire w103036;
	repeater #(1, 1'b0, 0, 0) c103036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103036));
	wire w105036;
	torch #(1'b0) c105036 (.i_clk(tick), .i_in(), .o_out(w105036));
	wire w121036;

	wire w122036;

	wire w135036;

	wire w159036;

	wire w172036;

	wire w173036;

	wire w120037;

	wire w129037;

	wire w165037;

	wire w174037;

	wire w73038;
	repeater #(1, 1'b0, 0, 0) c73038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73038));
	wire w107038;
	repeater #(1, 1'b0, 0, 0) c107038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107038));
	wire w123038;

	wire w153038;
	assign outputs[79] = ();
	wire w171038;

	wire w70040;
	torch #(1'b1) c70040 (.i_clk(tick), .i_in(), .o_out(w70040));
	wire w104040;
	torch #(1'b1) c104040 (.i_clk(tick), .i_in(), .o_out(w104040));
	wire w186040;

	wire w190040;

	wire w194040;

	wire w198040;

	wire w202040;

	wire w206040;

	wire w2041;

	wire w69043;
	repeater #(2, 1'b0, 0, 0) c69043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69043));
	wire w103043;
	repeater #(2, 1'b0, 0, 0) c103043 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103043));
	wire w49047;
	torch #(1'b0) c49047 (.i_clk(tick), .i_in(), .o_out(w49047));
	wire w50047;
	torch #(1'b0) c50047 (.i_clk(tick), .i_in(), .o_out(w50047));
	wire w57047;
	torch #(1'b0) c57047 (.i_clk(tick), .i_in(), .o_out(w57047));
	wire w58047;
	torch #(1'b0) c58047 (.i_clk(tick), .i_in(), .o_out(w58047));
	wire w65047;
	torch #(1'b0) c65047 (.i_clk(tick), .i_in(), .o_out(w65047));
	wire w66047;
	torch #(1'b0) c66047 (.i_clk(tick), .i_in(), .o_out(w66047));
	wire w73047;
	torch #(1'b0) c73047 (.i_clk(tick), .i_in(), .o_out(w73047));
	wire w74047;
	torch #(1'b0) c74047 (.i_clk(tick), .i_in(), .o_out(w74047));
	wire w83047;
	torch #(1'b0) c83047 (.i_clk(tick), .i_in(), .o_out(w83047));
	wire w84047;
	torch #(1'b0) c84047 (.i_clk(tick), .i_in(), .o_out(w84047));
	wire w91047;
	torch #(1'b0) c91047 (.i_clk(tick), .i_in(), .o_out(w91047));
	wire w92047;
	torch #(1'b0) c92047 (.i_clk(tick), .i_in(), .o_out(w92047));
	wire w99047;
	torch #(1'b0) c99047 (.i_clk(tick), .i_in(), .o_out(w99047));
	wire w100047;
	torch #(1'b0) c100047 (.i_clk(tick), .i_in(), .o_out(w100047));
	wire w107047;
	torch #(1'b0) c107047 (.i_clk(tick), .i_in(), .o_out(w107047));
	wire w108047;
	torch #(1'b0) c108047 (.i_clk(tick), .i_in(), .o_out(w108047));
	wire w186051;
	torch #(1'b0) c186051 (.i_clk(tick), .i_in(), .o_out(w186051));
	wire w190051;
	torch #(1'b0) c190051 (.i_clk(tick), .i_in(), .o_out(w190051));
	wire w194051;
	torch #(1'b0) c194051 (.i_clk(tick), .i_in(), .o_out(w194051));
	wire w198051;
	torch #(1'b0) c198051 (.i_clk(tick), .i_in(), .o_out(w198051));
	wire w202051;
	torch #(1'b0) c202051 (.i_clk(tick), .i_in(), .o_out(w202051));
	wire w206051;
	torch #(1'b0) c206051 (.i_clk(tick), .i_in(), .o_out(w206051));
	wire w2052;
	torch #(1'b0) c2052 (.i_clk(tick), .i_in(), .o_out(w2052));
	wire w94054;
	repeater #(1, 1'b0, 0, 0) c94054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94054));
	wire w186056;

	wire w190056;

	wire w194056;

	wire w198056;

	wire w202056;

	wire w206056;

	wire w2057;

	wire w140060;

	wire w158060;

	wire w186067;
	torch #(1'b0) c186067 (.i_clk(tick), .i_in(), .o_out(w186067));
	wire w190067;
	torch #(1'b0) c190067 (.i_clk(tick), .i_in(), .o_out(w190067));
	wire w194067;
	torch #(1'b0) c194067 (.i_clk(tick), .i_in(), .o_out(w194067));
	wire w198067;
	torch #(1'b0) c198067 (.i_clk(tick), .i_in(), .o_out(w198067));
	wire w202067;
	torch #(1'b0) c202067 (.i_clk(tick), .i_in(), .o_out(w202067));
	wire w206067;
	torch #(1'b0) c206067 (.i_clk(tick), .i_in(), .o_out(w206067));
	wire w2068;
	torch #(1'b0) c2068 (.i_clk(tick), .i_in(), .o_out(w2068));
	wire w186072;

	wire w190072;

	wire w194072;

	wire w198072;

	wire w202072;

	wire w206072;

	wire w2073;

	wire w186083;
	torch #(1'b0) c186083 (.i_clk(tick), .i_in(), .o_out(w186083));
	wire w190083;
	torch #(1'b0) c190083 (.i_clk(tick), .i_in(), .o_out(w190083));
	wire w194083;
	torch #(1'b0) c194083 (.i_clk(tick), .i_in(), .o_out(w194083));
	wire w198083;
	torch #(1'b0) c198083 (.i_clk(tick), .i_in(), .o_out(w198083));
	wire w202083;
	torch #(1'b0) c202083 (.i_clk(tick), .i_in(), .o_out(w202083));
	wire w206083;
	torch #(1'b0) c206083 (.i_clk(tick), .i_in(), .o_out(w206083));
	wire w2084;
	torch #(1'b0) c2084 (.i_clk(tick), .i_in(), .o_out(w2084));
	wire w184086;
	assign outputs[80] = ();
	wire w186086;
	assign outputs[81] = ();
	wire w188086;
	assign outputs[82] = ();
	wire w190086;
	assign outputs[83] = ();
	wire w192086;
	assign outputs[84] = ();
	wire w194086;
	assign outputs[85] = ();
	wire w196086;
	assign outputs[86] = ();
	wire w198086;
	assign outputs[87] = ();
	wire w200086;
	assign outputs[88] = ();
	wire w202086;
	assign outputs[89] = ();
	wire w204086;
	assign outputs[90] = ();
	wire w206086;
	assign outputs[91] = ();
	wire w0087;
	assign outputs[92] = ();
	wire w2087;
	assign outputs[93] = ();
	wire w184087;
	repeater #(1, 1'b0, 0, 0) c184087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184087));
	wire w186087;
	repeater #(1, 1'b0, 0, 0) c186087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186087));
	wire w188087;
	repeater #(1, 1'b0, 0, 0) c188087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188087));
	wire w190087;
	repeater #(1, 1'b0, 0, 0) c190087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190087));
	wire w192087;
	repeater #(1, 1'b0, 0, 0) c192087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192087));
	wire w194087;
	repeater #(1, 1'b0, 0, 0) c194087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194087));
	wire w196087;
	repeater #(1, 1'b0, 0, 0) c196087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196087));
	wire w198087;
	repeater #(1, 1'b0, 0, 0) c198087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198087));
	wire w200087;
	repeater #(1, 1'b0, 0, 0) c200087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200087));
	wire w202087;
	repeater #(1, 1'b0, 0, 0) c202087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202087));
	wire w204087;
	repeater #(1, 1'b0, 0, 0) c204087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w204087));
	wire w206087;
	repeater #(1, 1'b0, 0, 0) c206087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206087));
	wire w0088;
	repeater #(1, 1'b0, 0, 0) c0088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0088));
	wire w2088;
	repeater #(1, 1'b0, 0, 0) c2088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2088));
	wire w185094;
	repeater #(2, 1'b1, 0, 0) c185094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w185094));
	wire w189094;
	repeater #(2, 1'b1, 0, 0) c189094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w189094));
	wire w193094;
	repeater #(2, 1'b1, 0, 0) c193094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193094));
	wire w197094;
	repeater #(2, 1'b1, 0, 0) c197094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197094));
	wire w201094;
	repeater #(2, 1'b1, 0, 0) c201094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w201094));
	wire w205094;
	repeater #(2, 1'b1, 0, 0) c205094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w205094));
	wire w1095;
	repeater #(2, 1'b1, 0, 0) c1095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1095));
	wire w183099;
	repeater #(1, 1'b1, 0, 0) c183099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183099));
	wire w187099;
	repeater #(1, 1'b1, 0, 0) c187099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187099));
	wire w191099;
	repeater #(1, 1'b1, 0, 0) c191099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191099));
	wire w195099;
	repeater #(1, 1'b1, 0, 0) c195099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195099));
	wire w199099;
	repeater #(1, 1'b1, 0, 0) c199099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199099));
	wire w203099;
	repeater #(1, 1'b1, 0, 0) c203099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203099));
	wire w207099;
	repeater #(1, 1'b1, 0, 0) c207099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207099));
	wire w1850100;

	wire w1890100;

	wire w1930100;

	wire w1970100;

	wire w2010100;

	wire w2050100;

	wire w10101;

	wire w1840101;

	wire w1880101;

	wire w1920101;

	wire w1960101;

	wire w2000101;

	wire w2040101;

	wire w00102;

	wire w1850102;
	torch #(1'b1) c1850102 (.i_clk(tick), .i_in(), .o_out(w1850102));
	wire w1890102;
	torch #(1'b1) c1890102 (.i_clk(tick), .i_in(), .o_out(w1890102));
	wire w1930102;
	torch #(1'b1) c1930102 (.i_clk(tick), .i_in(), .o_out(w1930102));
	wire w1970102;
	torch #(1'b1) c1970102 (.i_clk(tick), .i_in(), .o_out(w1970102));
	wire w2010102;
	torch #(1'b1) c2010102 (.i_clk(tick), .i_in(), .o_out(w2010102));
	wire w2050102;
	torch #(1'b1) c2050102 (.i_clk(tick), .i_in(), .o_out(w2050102));
	wire w10103;
	torch #(1'b1) c10103 (.i_clk(tick), .i_in(), .o_out(w10103));
	wire w1830103;
	repeater #(1, 1'b1, 0, 0) c1830103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830103));
	wire w1870103;
	repeater #(1, 1'b1, 0, 0) c1870103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870103));
	wire w1910103;
	repeater #(1, 1'b1, 0, 0) c1910103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910103));
	wire w1950103;
	repeater #(1, 1'b1, 0, 0) c1950103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1950103));
	wire w1990103;
	repeater #(1, 1'b1, 0, 0) c1990103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990103));
	wire w2030103;
	repeater #(1, 1'b1, 0, 0) c2030103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030103));
	wire w2070103;
	repeater #(1, 1'b1, 0, 0) c2070103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070103));
	wire w40115;
	torch #(1'b1) c40115 (.i_clk(tick), .i_in(), .o_out(w40115));
	wire w1860115;
	torch #(1'b1) c1860115 (.i_clk(tick), .i_in(), .o_out(w1860115));
	wire w1900115;
	torch #(1'b1) c1900115 (.i_clk(tick), .i_in(), .o_out(w1900115));
	wire w1940115;
	torch #(1'b1) c1940115 (.i_clk(tick), .i_in(), .o_out(w1940115));
	wire w1980115;
	torch #(1'b1) c1980115 (.i_clk(tick), .i_in(), .o_out(w1980115));
	wire w2020115;
	torch #(1'b1) c2020115 (.i_clk(tick), .i_in(), .o_out(w2020115));
	wire w2060115;
	torch #(1'b1) c2060115 (.i_clk(tick), .i_in(), .o_out(w2060115));
	wire w20116;
	torch #(1'b1) c20116 (.i_clk(tick), .i_in(), .o_out(w20116));
	wire w20162;

	wire w00164;

	wire w2060165;

	wire w2040167;

	wire w2020169;

	wire w600174;
	repeater #(2, 1'b1, 0, 0) c600174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600174));
	wire w940174;
	repeater #(2, 1'b1, 0, 0) c940174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w940174));
	wire w1850175;
	torch #(1'b1) c1850175 (.i_clk(tick), .i_in(), .o_out(w1850175));
	wire w1890175;
	torch #(1'b1) c1890175 (.i_clk(tick), .i_in(), .o_out(w1890175));
	wire w1930175;
	torch #(1'b1) c1930175 (.i_clk(tick), .i_in(), .o_out(w1930175));
	wire w1970175;
	torch #(1'b1) c1970175 (.i_clk(tick), .i_in(), .o_out(w1970175));
	wire w2010175;
	torch #(1'b1) c2010175 (.i_clk(tick), .i_in(), .o_out(w2010175));
	wire w2050175;
	torch #(1'b1) c2050175 (.i_clk(tick), .i_in(), .o_out(w2050175));
	wire w10176;
	torch #(1'b1) c10176 (.i_clk(tick), .i_in(), .o_out(w10176));
	wire w520176;
	torch #(1'b1) c520176 (.i_clk(tick), .i_in(), .o_out(w520176));
	wire w620176;
	repeater #(1, 1'b1, 0, 0) c620176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620176));
	wire w860176;
	torch #(1'b1) c860176 (.i_clk(tick), .i_in(), .o_out(w860176));
	wire w960176;
	repeater #(1, 1'b1, 0, 0) c960176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w960176));
	wire w1860178;
	repeater #(2, 1'b0, 0, 0) c1860178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1860178));
	wire w1900178;
	repeater #(2, 1'b0, 0, 0) c1900178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1900178));
	wire w1940178;
	repeater #(2, 1'b0, 0, 0) c1940178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1940178));
	wire w1980178;
	repeater #(2, 1'b0, 0, 0) c1980178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980178));
	wire w2020178;
	repeater #(1, 1'b0, 0, 0) c2020178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020178));
	wire w2060178;
	repeater #(1, 1'b0, 0, 0) c2060178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060178));
	wire w210;
	repeater #(1, 1'b0, 0, 0) c210 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w210));
	wire w19910;
	repeater #(1, 1'b0, 0, 0) c19910 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19910));
	wire w311;
	repeater #(1, 1'b0, 0, 0) c311 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w311));
	wire w6211;
	repeater #(1, 1'b1, 0, 0) c6211 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6211));
	wire w9611;
	repeater #(1, 1'b1, 0, 0) c9611 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9611));
	wire w5112;

	wire w8512;

	wire w6114;

	wire w6214;

	wire w9514;

	wire w9614;

	wire w18815;
	repeater #(1, 1'b0, 0, 0) c18815 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18815));
	wire w016;
	repeater #(1, 1'b0, 0, 0) c016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w016));
	wire w5416;

	wire w8816;

	wire w6017;

	wire w6117;

	wire w9417;

	wire w9517;

	wire w4618;

	wire w8018;

	wire w12318;
	repeater #(2, 1'b1, 0, 0) c12318 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12318));
	wire w12518;
	repeater #(1, 1'b1, 0, 0) c12518 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12518));
	wire w12718;
	repeater #(2, 1'b1, 0, 0) c12718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12718));
	wire w12918;
	repeater #(1, 1'b0, 0, 0) c12918 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12918));
	wire w13118;
	repeater #(2, 1'b1, 0, 0) c13118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13118));
	wire w13318;
	repeater #(1, 1'b1, 0, 0) c13318 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13318));
	wire w13518;
	repeater #(2, 1'b1, 0, 0) c13518 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13518));
	wire w13718;
	repeater #(1, 1'b1, 0, 0) c13718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13718));
	wire w15718;
	repeater #(1, 1'b1, 0, 0) c15718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15718));
	wire w15918;
	repeater #(2, 1'b1, 0, 0) c15918 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15918));
	wire w16118;
	repeater #(1, 1'b1, 0, 0) c16118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16118));
	wire w16318;
	repeater #(2, 1'b1, 0, 0) c16318 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16318));
	wire w16518;
	repeater #(1, 1'b1, 0, 0) c16518 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16518));
	wire w16718;
	repeater #(2, 1'b1, 0, 0) c16718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16718));
	wire w16918;
	repeater #(1, 1'b1, 0, 0) c16918 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16918));
	wire w17118;
	repeater #(2, 1'b1, 0, 0) c17118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17118));
	wire w18318;
	repeater #(2, 1'b0, 0, 0) c18318 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18318));
	wire w47110;
	repeater #(1, 1'b1, 0, 0) c47110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47110));
	wire w51110;
	repeater #(1, 1'b1, 0, 0) c51110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51110));
	wire w55110;
	repeater #(1, 1'b1, 0, 0) c55110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55110));
	wire w59110;
	repeater #(1, 1'b1, 0, 0) c59110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59110));
	wire w63110;
	repeater #(1, 1'b1, 0, 0) c63110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63110));
	wire w67110;
	repeater #(1, 1'b1, 0, 0) c67110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67110));
	wire w71110;
	repeater #(1, 1'b1, 0, 0) c71110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71110));
	wire w81110;
	repeater #(1, 1'b1, 0, 0) c81110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81110));
	wire w85110;
	repeater #(1, 1'b1, 0, 0) c85110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85110));
	wire w89110;
	repeater #(1, 1'b1, 0, 0) c89110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89110));
	wire w93110;
	repeater #(1, 1'b1, 0, 0) c93110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93110));
	wire w97110;
	repeater #(1, 1'b1, 0, 0) c97110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97110));
	wire w101110;
	repeater #(1, 1'b1, 0, 0) c101110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101110));
	wire w105110;
	repeater #(1, 1'b1, 0, 0) c105110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105110));
	wire w132110;

	wire w162110;

	wire w124111;

	wire w128111;

	wire w131111;

	wire w133111;

	wire w136111;

	wire w158111;

	wire w161111;

	wire w163111;

	wire w166111;

	wire w170111;

	wire w123112;

	wire w125112;

	wire w127112;

	wire w129112;

	wire w132112;

	wire w135112;

	wire w137112;

	wire w157112;

	wire w159112;

	wire w162112;

	wire w165112;

	wire w167112;

	wire w169112;

	wire w171112;

	wire w128113;

	wire w145113;
	repeater #(1, 1'b1, 0, 0) c145113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145113));
	wire w166113;

	wire w184113;
	torch #(1'b1) c184113 (.i_clk(tick), .i_in(), .o_out(w184113));
	wire w188113;
	torch #(1'b1) c188113 (.i_clk(tick), .i_in(), .o_out(w188113));
	wire w192113;
	torch #(1'b1) c192113 (.i_clk(tick), .i_in(), .o_out(w192113));
	wire w196113;
	torch #(1'b1) c196113 (.i_clk(tick), .i_in(), .o_out(w196113));
	wire w200113;
	torch #(1'b1) c200113 (.i_clk(tick), .i_in(), .o_out(w200113));
	wire w204113;
	torch #(1'b1) c204113 (.i_clk(tick), .i_in(), .o_out(w204113));
	wire w0114;
	torch #(1'b1) c0114 (.i_clk(tick), .i_in(), .o_out(w0114));
	wire w124114;

	wire w128114;

	wire w129114;

	wire w133114;

	wire w135114;

	wire w137114;

	wire w157114;

	wire w159114;

	wire w161114;

	wire w165114;

	wire w166114;

	wire w170114;

	wire w125116;

	wire w127116;

	wire w129116;

	wire w165116;

	wire w167116;

	wire w169116;

	wire w59121;
	repeater #(1, 1'b1, 0, 0) c59121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w59121));
	wire w93121;
	repeater #(1, 1'b1, 0, 0) c93121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w93121));
	wire w188121;
	repeater #(1, 1'b0, 0, 0) c188121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188121));
	wire w0122;
	repeater #(1, 1'b0, 0, 0) c0122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0122));
	wire w70122;

	wire w104122;

	wire w59124;

	wire w73124;

	wire w93124;

	wire w107124;

	wire w183124;
	repeater #(2, 1'b0, 0, 0) c183124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183124));
	wire w59128;

	wire w60128;

	wire w73128;

	wire w93128;

	wire w94128;

	wire w107128;

	wire w184129;
	torch #(1'b1) c184129 (.i_clk(tick), .i_in(), .o_out(w184129));
	wire w188129;
	torch #(1'b1) c188129 (.i_clk(tick), .i_in(), .o_out(w188129));
	wire w192129;
	torch #(1'b1) c192129 (.i_clk(tick), .i_in(), .o_out(w192129));
	wire w196129;
	torch #(1'b1) c196129 (.i_clk(tick), .i_in(), .o_out(w196129));
	wire w200129;
	torch #(1'b1) c200129 (.i_clk(tick), .i_in(), .o_out(w200129));
	wire w204129;
	torch #(1'b1) c204129 (.i_clk(tick), .i_in(), .o_out(w204129));
	wire w0130;
	torch #(1'b1) c0130 (.i_clk(tick), .i_in(), .o_out(w0130));
	wire w70130;
	torch #(1'b1) c70130 (.i_clk(tick), .i_in(), .o_out(w70130));
	wire w71130;

	wire w104130;
	torch #(1'b1) c104130 (.i_clk(tick), .i_in(), .o_out(w104130));
	wire w105130;

	wire w120130;
	repeater #(2, 1'b0, 0, 0) c120130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120130));
	wire w147130;

	wire w174130;
	repeater #(2, 1'b0, 0, 0) c174130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174130));
	wire w71131;

	wire w73131;

	wire w105131;

	wire w107131;

	wire w118131;

	wire w119131;

	wire w125131;
	repeater #(1, 1'b1, 0, 0) c125131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125131));
	wire w126131;
	repeater #(2, 1'b1, 0, 0) c126131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126131));
	wire w148131;

	wire w168131;
	repeater #(2, 1'b1, 0, 0) c168131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168131));
	wire w169131;
	repeater #(1, 1'b1, 0, 0) c169131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169131));
	wire w175131;

	wire w176131;

	wire w122132;
	repeater #(2, 1'b1, 0, 0) c122132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122132));
	wire w123132;
	repeater #(2, 1'b1, 0, 0) c123132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123132));
	wire w125132;

	wire w148132;
	repeater #(1, 1'b1, 0, 0) c148132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148132));
	wire w169132;

	wire w171132;
	repeater #(2, 1'b1, 0, 0) c171132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171132));
	wire w172132;
	repeater #(2, 1'b1, 0, 0) c172132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172132));
	wire w73133;

	wire w74133;

	wire w75133;

	wire w107133;

	wire w108133;

	wire w109133;

	wire w123133;

	wire w125133;
	repeater #(1, 1'b1, 0, 0) c125133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125133));
	wire w136133;

	wire w137133;

	wire w157133;

	wire w158133;

	wire w169133;
	repeater #(1, 1'b1, 0, 0) c169133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169133));
	wire w171133;

	wire w68134;

	wire w69134;

	wire w75134;

	wire w102134;

	wire w103134;

	wire w109134;

	wire w119134;

	wire w123134;

	wire w147134;

	wire w148134;

	wire w171134;

	wire w175134;

	wire w119135;

	wire w121135;
	repeater #(1, 1'b0, 0, 0) c121135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121135));
	wire w126135;

	wire w130135;

	wire w136135;
	repeater #(1, 1'b0, 0, 0) c136135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136135));
	wire w158135;
	repeater #(1, 1'b0, 0, 0) c158135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158135));
	wire w164135;

	wire w168135;

	wire w173135;
	repeater #(1, 1'b1, 0, 0) c173135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173135));
	wire w175135;

	wire w73136;
	repeater #(1, 1'b0, 0, 0) c73136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73136));
	wire w75136;
	torch #(1'b0) c75136 (.i_clk(tick), .i_in(), .o_out(w75136));
	wire w107136;
	repeater #(1, 1'b0, 0, 0) c107136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107136));
	wire w109136;
	torch #(1'b0) c109136 (.i_clk(tick), .i_in(), .o_out(w109136));
	wire w126136;

	wire w128136;
	repeater #(1, 1'b0, 0, 0) c128136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128136));
	wire w129136;

	wire w136136;

	wire w153136;

	wire w158136;

	wire w165136;

	wire w166136;
	repeater #(1, 1'b1, 0, 0) c166136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166136));
	wire w168136;

	wire w122137;

	wire w137137;

	wire w141137;
	repeater #(1, 1'b0, 0, 0) c141137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141137));
	wire w154137;
	repeater #(2, 1'b0, 0, 0) c154137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154137));
	wire w157137;

	wire w172137;

	wire w188137;
	repeater #(1, 1'b0, 0, 0) c188137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188137));
	wire w0138;
	repeater #(1, 1'b0, 0, 0) c0138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0138));
	wire w119138;

	wire w120138;
	repeater #(1, 1'b1, 0, 0) c120138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120138));
	wire w127138;
	repeater #(2, 1'b1, 0, 0) c127138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127138));
	wire w140138;
	assign outputs[94] = ();
	wire w167138;
	repeater #(2, 1'b1, 0, 0) c167138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167138));
	wire w174138;
	repeater #(1, 1'b0, 0, 0) c174138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174138));
	wire w175138;

	wire w74140;
	torch #(1'b1) c74140 (.i_clk(tick), .i_in(), .o_out(w74140));
	wire w108140;
	torch #(1'b1) c108140 (.i_clk(tick), .i_in(), .o_out(w108140));
	wire w183140;
	repeater #(2, 1'b0, 0, 0) c183140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183140));
	wire w73143;
	repeater #(2, 1'b0, 0, 0) c73143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73143));
	wire w107143;
	repeater #(2, 1'b0, 0, 0) c107143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107143));
	wire w184145;
	torch #(1'b1) c184145 (.i_clk(tick), .i_in(), .o_out(w184145));
	wire w188145;
	torch #(1'b1) c188145 (.i_clk(tick), .i_in(), .o_out(w188145));
	wire w192145;
	torch #(1'b1) c192145 (.i_clk(tick), .i_in(), .o_out(w192145));
	wire w196145;
	torch #(1'b1) c196145 (.i_clk(tick), .i_in(), .o_out(w196145));
	wire w200145;
	torch #(1'b1) c200145 (.i_clk(tick), .i_in(), .o_out(w200145));
	wire w204145;
	torch #(1'b1) c204145 (.i_clk(tick), .i_in(), .o_out(w204145));
	wire w0146;
	torch #(1'b1) c0146 (.i_clk(tick), .i_in(), .o_out(w0146));
	wire w188153;
	repeater #(1, 1'b0, 0, 0) c188153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188153));
	wire w0154;
	repeater #(1, 1'b0, 0, 0) c0154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0154));
	wire w63156;
	repeater #(1, 1'b0, 0, 0) c63156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63156));
	wire w183156;
	repeater #(2, 1'b0, 0, 0) c183156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183156));
	wire w148161;
	repeater #(1, 1'b0, 0, 0) c148161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148161));
	wire w151161;
	repeater #(2, 1'b0, 0, 0) c151161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151161));
	wire w184161;
	torch #(1'b1) c184161 (.i_clk(tick), .i_in(), .o_out(w184161));
	wire w188161;
	torch #(1'b1) c188161 (.i_clk(tick), .i_in(), .o_out(w188161));
	wire w192161;
	torch #(1'b1) c192161 (.i_clk(tick), .i_in(), .o_out(w192161));
	wire w196161;
	torch #(1'b1) c196161 (.i_clk(tick), .i_in(), .o_out(w196161));
	wire w200161;
	torch #(1'b1) c200161 (.i_clk(tick), .i_in(), .o_out(w200161));
	wire w204161;
	torch #(1'b1) c204161 (.i_clk(tick), .i_in(), .o_out(w204161));
	wire w0162;
	torch #(1'b1) c0162 (.i_clk(tick), .i_in(), .o_out(w0162));
	wire w143162;
	repeater #(1, 1'b0, 0, 0) c143162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143162));
	wire w156162;
	repeater #(2, 1'b0, 0, 0) c156162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156162));
	wire w142163;
	assign outputs[95] = ();
	wire w145163;

	wire w154163;

	wire w145164;

	wire w154164;

	wire w143165;
	repeater #(1, 1'b0, 0, 0) c143165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143165));
	wire w156165;
	repeater #(1, 1'b0, 0, 0) c156165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156165));
	wire w188169;
	repeater #(1, 1'b0, 0, 0) c188169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188169));
	wire w0170;
	repeater #(1, 1'b0, 0, 0) c0170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0170));
	wire w183172;
	repeater #(2, 1'b0, 0, 0) c183172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183172));
	wire w184177;
	torch #(1'b1) c184177 (.i_clk(tick), .i_in(), .o_out(w184177));
	wire w188177;
	torch #(1'b1) c188177 (.i_clk(tick), .i_in(), .o_out(w188177));
	wire w192177;
	torch #(1'b1) c192177 (.i_clk(tick), .i_in(), .o_out(w192177));
	wire w196177;
	torch #(1'b1) c196177 (.i_clk(tick), .i_in(), .o_out(w196177));
	wire w200177;
	torch #(1'b1) c200177 (.i_clk(tick), .i_in(), .o_out(w200177));
	wire w204177;
	torch #(1'b1) c204177 (.i_clk(tick), .i_in(), .o_out(w204177));
	wire w0178;
	torch #(1'b1) c0178 (.i_clk(tick), .i_in(), .o_out(w0178));
	wire w183190;
	repeater #(1, 1'b0, 0, 0) c183190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183190));
	wire w185190;
	torch #(1'b1) c185190 (.i_clk(tick), .i_in(), .o_out(w185190));
	wire w187190;
	repeater #(1, 1'b0, 0, 0) c187190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187190));
	wire w189190;
	torch #(1'b1) c189190 (.i_clk(tick), .i_in(), .o_out(w189190));
	wire w191190;
	repeater #(1, 1'b0, 0, 0) c191190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191190));
	wire w193190;
	torch #(1'b1) c193190 (.i_clk(tick), .i_in(), .o_out(w193190));
	wire w195190;
	repeater #(1, 1'b0, 0, 0) c195190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w195190));
	wire w197190;
	torch #(1'b1) c197190 (.i_clk(tick), .i_in(), .o_out(w197190));
	wire w199190;
	repeater #(1, 1'b0, 0, 0) c199190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199190));
	wire w201190;
	torch #(1'b1) c201190 (.i_clk(tick), .i_in(), .o_out(w201190));
	wire w203190;
	repeater #(1, 1'b0, 0, 0) c203190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w203190));
	wire w205190;
	torch #(1'b1) c205190 (.i_clk(tick), .i_in(), .o_out(w205190));
	wire w207190;
	repeater #(1, 1'b0, 0, 0) c207190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207190));
	wire w1191;
	torch #(1'b1) c1191 (.i_clk(tick), .i_in(), .o_out(w1191));
	wire w185194;
	torch #(1'b1) c185194 (.i_clk(tick), .i_in(), .o_out(w185194));
	wire w189194;
	torch #(1'b1) c189194 (.i_clk(tick), .i_in(), .o_out(w189194));
	wire w193194;
	torch #(1'b1) c193194 (.i_clk(tick), .i_in(), .o_out(w193194));
	wire w197194;
	torch #(1'b1) c197194 (.i_clk(tick), .i_in(), .o_out(w197194));
	wire w201194;
	torch #(1'b1) c201194 (.i_clk(tick), .i_in(), .o_out(w201194));
	wire w205194;
	torch #(1'b1) c205194 (.i_clk(tick), .i_in(), .o_out(w205194));
	wire w1195;
	torch #(1'b1) c1195 (.i_clk(tick), .i_in(), .o_out(w1195));
	wire w1841102;
	torch #(1'b1) c1841102 (.i_clk(tick), .i_in(), .o_out(w1841102));
	wire w1881102;
	torch #(1'b1) c1881102 (.i_clk(tick), .i_in(), .o_out(w1881102));
	wire w1921102;
	torch #(1'b1) c1921102 (.i_clk(tick), .i_in(), .o_out(w1921102));
	wire w1961102;
	torch #(1'b1) c1961102 (.i_clk(tick), .i_in(), .o_out(w1961102));
	wire w2001102;
	torch #(1'b1) c2001102 (.i_clk(tick), .i_in(), .o_out(w2001102));
	wire w2041102;
	torch #(1'b1) c2041102 (.i_clk(tick), .i_in(), .o_out(w2041102));
	wire w01103;
	torch #(1'b1) c01103 (.i_clk(tick), .i_in(), .o_out(w01103));
	wire w1911116;
	repeater #(1, 1'b0, 0, 0) c1911116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911116));
	wire w1991116;
	repeater #(1, 1'b0, 0, 0) c1991116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991116));
	wire w2071116;
	repeater #(1, 1'b0, 0, 0) c2071116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071116));
	wire w1931118;
	repeater #(1, 1'b0, 0, 0) c1931118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1931118));
	wire w1991118;
	repeater #(1, 1'b0, 0, 0) c1991118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991118));
	wire w11119;
	repeater #(1, 1'b0, 0, 0) c11119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11119));
	wire w2011120;
	repeater #(1, 1'b0, 0, 0) c2011120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2011120));
	wire w2051120;
	repeater #(1, 1'b0, 0, 0) c2051120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2051120));
	wire w11121;
	repeater #(1, 1'b0, 0, 0) c11121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11121));
	wire w1851135;
	repeater #(1, 1'b0, 0, 0) c1851135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1851135));
	wire w1891135;
	repeater #(1, 1'b0, 0, 0) c1891135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1891135));
	wire w1931135;
	repeater #(1, 1'b0, 0, 0) c1931135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1931135));
	wire w1971135;
	repeater #(1, 1'b0, 0, 0) c1971135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1971135));
	wire w2011135;
	repeater #(1, 1'b0, 0, 0) c2011135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2011135));
	wire w2051135;
	repeater #(1, 1'b0, 0, 0) c2051135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2051135));
	wire w11136;
	repeater #(1, 1'b0, 0, 0) c11136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11136));
	wire w16902;
	torch #(1'b1) c16902 (.i_clk(tick), .i_in(), .o_out(w16902));
	wire w17302;
	torch #(1'b1) c17302 (.i_clk(tick), .i_in(), .o_out(w17302));
	wire w17702;
	torch #(1'b1) c17702 (.i_clk(tick), .i_in(), .o_out(w17702));
	wire w18102;
	torch #(1'b1) c18102 (.i_clk(tick), .i_in(), .o_out(w18102));
	wire w18502;
	torch #(1'b1) c18502 (.i_clk(tick), .i_in(), .o_out(w18502));
	wire w18902;
	torch #(1'b1) c18902 (.i_clk(tick), .i_in(), .o_out(w18902));
	wire w19302;
	torch #(1'b1) c19302 (.i_clk(tick), .i_in(), .o_out(w19302));
	wire w18005;
	repeater #(1, 1'b1, 0, 0) c18005 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18005));
	wire w18205;
	repeater #(1, 1'b1, 0, 0) c18205 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18205));
	wire w18405;
	repeater #(1, 1'b1, 0, 0) c18405 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18405));
	wire w18605;
	repeater #(1, 1'b1, 0, 0) c18605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18605));
	wire w18805;
	repeater #(1, 1'b1, 0, 0) c18805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18805));
	wire w19005;
	repeater #(1, 1'b1, 0, 0) c19005 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19005));
	wire w19205;
	repeater #(1, 1'b1, 0, 0) c19205 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19205));
	wire w19405;
	repeater #(1, 1'b1, 0, 0) c19405 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19405));
	wire w17807;
	repeater #(1, 1'b1, 0, 0) c17807 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17807));
	wire w17609;
	repeater #(1, 1'b1, 0, 0) c17609 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17609));
	wire w174011;
	repeater #(1, 1'b1, 0, 0) c174011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174011));
	wire w172013;
	repeater #(1, 1'b1, 0, 0) c172013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172013));
	wire w170015;
	repeater #(1, 1'b1, 0, 0) c170015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170015));
	wire w114016;
	repeater #(1, 1'b1, 0, 0) c114016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114016));
	wire w168017;
	repeater #(1, 1'b1, 0, 0) c168017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168017));
	wire w58023;
	torch #(1'b1) c58023 (.i_clk(tick), .i_in(), .o_out(w58023));
	wire w92023;
	repeater #(1, 1'b1, 0, 0) c92023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92023));
	wire w126023;
	torch #(1'b1) c126023 (.i_clk(tick), .i_in(), .o_out(w126023));
	wire w160023;
	repeater #(1, 1'b1, 0, 0) c160023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160023));
	wire w56025;
	repeater #(1, 1'b1, 0, 0) c56025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56025));
	wire w90025;
	repeater #(1, 1'b1, 0, 0) c90025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90025));
	wire w105025;
	repeater #(1, 1'b1, 0, 0) c105025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105025));
	wire w124025;
	repeater #(1, 1'b1, 0, 0) c124025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124025));
	wire w158025;
	repeater #(1, 1'b1, 0, 0) c158025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158025));
	wire w194026;
	repeater #(1, 1'b1, 0, 0) c194026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194026));
	wire w54027;
	torch #(1'b1) c54027 (.i_clk(tick), .i_in(), .o_out(w54027));
	wire w88027;
	repeater #(1, 1'b1, 0, 0) c88027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88027));
	wire w122027;
	torch #(1'b1) c122027 (.i_clk(tick), .i_in(), .o_out(w122027));
	wire w156027;
	repeater #(1, 1'b1, 0, 0) c156027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156027));
	wire w192028;
	repeater #(1, 1'b1, 0, 0) c192028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192028));
	wire w52029;
	repeater #(1, 1'b1, 0, 0) c52029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52029));
	wire w86029;
	repeater #(1, 1'b1, 0, 0) c86029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86029));
	wire w120029;
	repeater #(1, 1'b1, 0, 0) c120029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120029));
	wire w154029;
	repeater #(1, 1'b1, 0, 0) c154029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154029));
	wire w190030;
	repeater #(1, 1'b1, 0, 0) c190030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190030));
	wire w50031;
	torch #(1'b1) c50031 (.i_clk(tick), .i_in(), .o_out(w50031));
	wire w84031;
	repeater #(1, 1'b1, 0, 0) c84031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84031));
	wire w118031;
	torch #(1'b1) c118031 (.i_clk(tick), .i_in(), .o_out(w118031));
	wire w152031;
	repeater #(1, 1'b1, 0, 0) c152031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152031));
	wire w188032;
	repeater #(1, 1'b1, 0, 0) c188032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188032));
	wire w48033;
	repeater #(1, 1'b1, 0, 0) c48033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48033));
	wire w82033;
	repeater #(1, 1'b1, 0, 0) c82033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82033));
	wire w116033;
	repeater #(1, 1'b1, 0, 0) c116033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116033));
	wire w150033;
	repeater #(1, 1'b1, 0, 0) c150033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150033));
	wire w32034;
	repeater #(1, 1'b1, 0, 0) c32034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32034));
	wire w34034;
	torch #(1'b1) c34034 (.i_clk(tick), .i_in(), .o_out(w34034));
	wire w36034;
	repeater #(1, 1'b1, 0, 0) c36034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36034));
	wire w38034;
	torch #(1'b1) c38034 (.i_clk(tick), .i_in(), .o_out(w38034));
	wire w40034;
	repeater #(1, 1'b1, 0, 0) c40034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40034));
	wire w42034;
	torch #(1'b1) c42034 (.i_clk(tick), .i_in(), .o_out(w42034));
	wire w44034;
	repeater #(1, 1'b1, 0, 0) c44034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44034));
	wire w46034;
	torch #(1'b1) c46034 (.i_clk(tick), .i_in(), .o_out(w46034));
	wire w66034;
	repeater #(1, 1'b1, 0, 0) c66034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66034));
	wire w68034;
	repeater #(1, 1'b1, 0, 0) c68034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68034));
	wire w70034;
	repeater #(1, 1'b1, 0, 0) c70034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70034));
	wire w72034;
	repeater #(1, 1'b1, 0, 0) c72034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72034));
	wire w74034;
	repeater #(1, 1'b1, 0, 0) c74034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74034));
	wire w76034;
	repeater #(1, 1'b1, 0, 0) c76034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76034));
	wire w78034;
	repeater #(1, 1'b1, 0, 0) c78034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78034));
	wire w80034;
	repeater #(1, 1'b1, 0, 0) c80034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80034));
	wire w97034;
	assign w97034 = inputs[20];
	wire w102034;
	torch #(1'b1) c102034 (.i_clk(tick), .i_in(), .o_out(w102034));
	wire w106034;
	torch #(1'b1) c106034 (.i_clk(tick), .i_in(), .o_out(w106034));
	wire w110034;
	torch #(1'b1) c110034 (.i_clk(tick), .i_in(), .o_out(w110034));
	wire w114034;
	torch #(1'b1) c114034 (.i_clk(tick), .i_in(), .o_out(w114034));
	wire w134034;
	repeater #(1, 1'b1, 0, 0) c134034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134034));
	wire w136034;
	repeater #(1, 1'b1, 0, 0) c136034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136034));
	wire w138034;
	repeater #(1, 1'b1, 0, 0) c138034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138034));
	wire w140034;
	repeater #(1, 1'b1, 0, 0) c140034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140034));
	wire w142034;
	repeater #(1, 1'b1, 0, 0) c142034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142034));
	wire w144034;
	repeater #(1, 1'b1, 0, 0) c144034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144034));
	wire w146034;
	repeater #(1, 1'b1, 0, 0) c146034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146034));
	wire w148034;
	repeater #(1, 1'b1, 0, 0) c148034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148034));
	wire w186034;
	repeater #(1, 1'b1, 0, 0) c186034 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186034));
	wire w101035;
	repeater #(1, 1'b1, 0, 0) c101035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101035));
	wire w105035;
	repeater #(1, 1'b1, 0, 0) c105035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105035));
	wire w109035;
	repeater #(1, 1'b1, 0, 0) c109035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109035));
	wire w113035;
	repeater #(1, 1'b1, 0, 0) c113035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113035));
	wire w172035;
	repeater #(1, 1'b1, 0, 0) c172035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172035));
	wire w174035;
	repeater #(1, 1'b1, 0, 0) c174035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174035));
	wire w176035;
	repeater #(1, 1'b1, 0, 0) c176035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176035));
	wire w178035;
	repeater #(1, 1'b1, 0, 0) c178035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178035));
	wire w180035;
	repeater #(1, 1'b1, 0, 0) c180035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180035));
	wire w182035;
	repeater #(1, 1'b1, 0, 0) c182035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182035));
	wire w184035;
	repeater #(1, 1'b1, 0, 0) c184035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184035));
	wire w102037;
	torch #(1'b1) c102037 (.i_clk(tick), .i_in(), .o_out(w102037));
	wire w106037;
	torch #(1'b1) c106037 (.i_clk(tick), .i_in(), .o_out(w106037));
	wire w110037;
	torch #(1'b1) c110037 (.i_clk(tick), .i_in(), .o_out(w110037));
	wire w114037;
	torch #(1'b1) c114037 (.i_clk(tick), .i_in(), .o_out(w114037));
	wire w118037;
	torch #(1'b1) c118037 (.i_clk(tick), .i_in(), .o_out(w118037));
	wire w122037;
	torch #(1'b1) c122037 (.i_clk(tick), .i_in(), .o_out(w122037));
	wire w126037;
	torch #(1'b1) c126037 (.i_clk(tick), .i_in(), .o_out(w126037));
	wire w136037;
	torch #(1'b1) c136037 (.i_clk(tick), .i_in(), .o_out(w136037));
	wire w140037;
	torch #(1'b1) c140037 (.i_clk(tick), .i_in(), .o_out(w140037));
	wire w144037;
	torch #(1'b1) c144037 (.i_clk(tick), .i_in(), .o_out(w144037));
	wire w148037;
	torch #(1'b1) c148037 (.i_clk(tick), .i_in(), .o_out(w148037));
	wire w152037;
	torch #(1'b1) c152037 (.i_clk(tick), .i_in(), .o_out(w152037));
	wire w156037;
	torch #(1'b1) c156037 (.i_clk(tick), .i_in(), .o_out(w156037));
	wire w160037;
	torch #(1'b1) c160037 (.i_clk(tick), .i_in(), .o_out(w160037));
	wire w32038;
	repeater #(2, 1'b1, 0, 0) c32038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32038));
	wire w36038;
	repeater #(2, 1'b1, 0, 0) c36038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36038));
	wire w40038;
	repeater #(2, 1'b1, 0, 0) c40038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40038));
	wire w66038;
	repeater #(2, 1'b1, 0, 0) c66038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66038));
	wire w70038;
	repeater #(2, 1'b1, 0, 0) c70038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70038));
	wire w74038;
	repeater #(2, 1'b1, 0, 0) c74038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74038));
	wire w32040;
	torch #(1'b1) c32040 (.i_clk(tick), .i_in(), .o_out(w32040));
	wire w42040;
	repeater #(1, 1'b1, 0, 0) c42040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42040));
	wire w66040;
	torch #(1'b1) c66040 (.i_clk(tick), .i_in(), .o_out(w66040));
	wire w76040;
	repeater #(1, 1'b1, 0, 0) c76040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76040));
	wire w107041;
	torch #(1'b0) c107041 (.i_clk(tick), .i_in(), .o_out(w107041));
	wire w111041;
	torch #(1'b0) c111041 (.i_clk(tick), .i_in(), .o_out(w111041));
	wire w115041;
	torch #(1'b0) c115041 (.i_clk(tick), .i_in(), .o_out(w115041));
	wire w119041;
	torch #(1'b0) c119041 (.i_clk(tick), .i_in(), .o_out(w119041));
	wire w143041;
	torch #(1'b0) c143041 (.i_clk(tick), .i_in(), .o_out(w143041));
	wire w147041;
	torch #(1'b0) c147041 (.i_clk(tick), .i_in(), .o_out(w147041));
	wire w151041;
	torch #(1'b0) c151041 (.i_clk(tick), .i_in(), .o_out(w151041));
	wire w155041;
	torch #(1'b0) c155041 (.i_clk(tick), .i_in(), .o_out(w155041));
	wire w42044;
	repeater #(1, 1'b1, 0, 0) c42044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42044));
	wire w76044;
	repeater #(1, 1'b1, 0, 0) c76044 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76044));
	wire w31045;

	wire w65045;

	wire w170045;
	repeater #(1, 1'b1, 0, 0) c170045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170045));
	wire w174045;
	repeater #(1, 1'b1, 0, 0) c174045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174045));
	wire w178045;
	repeater #(1, 1'b1, 0, 0) c178045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178045));
	wire w182045;
	repeater #(1, 1'b1, 0, 0) c182045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182045));
	wire w186045;
	repeater #(1, 1'b1, 0, 0) c186045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186045));
	wire w190045;
	repeater #(1, 1'b1, 0, 0) c190045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190045));
	wire w194045;
	repeater #(1, 1'b1, 0, 0) c194045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194045));
	wire w42047;

	wire w76047;

	wire w34049;

	wire w68049;

	wire w172049;

	wire w197049;
	repeater #(2, 1'b0, 0, 0) c197049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197049));
	wire w40050;

	wire w41050;

	wire w74050;

	wire w75050;

	wire w192050;

	wire w176054;
	torch #(1'b1) c176054 (.i_clk(tick), .i_in(), .o_out(w176054));
	wire w180054;
	torch #(1'b1) c180054 (.i_clk(tick), .i_in(), .o_out(w180054));
	wire w184054;
	torch #(1'b1) c184054 (.i_clk(tick), .i_in(), .o_out(w184054));
	wire w188054;
	torch #(1'b1) c188054 (.i_clk(tick), .i_in(), .o_out(w188054));
	wire w31055;

	wire w32055;

	wire w35055;

	wire w36055;

	wire w39055;

	wire w40055;

	wire w43055;

	wire w44055;

	wire w47055;

	wire w48055;

	wire w51055;

	wire w52055;

	wire w55055;

	wire w56055;

	wire w65055;

	wire w66055;

	wire w69055;

	wire w70055;

	wire w73055;

	wire w74055;

	wire w77055;

	wire w78055;

	wire w81055;

	wire w82055;

	wire w85055;

	wire w86055;

	wire w89055;

	wire w90055;

	wire w130055;

	wire w32057;

	wire w36057;

	wire w40057;

	wire w44057;

	wire w48057;

	wire w52057;

	wire w56057;

	wire w66057;

	wire w70057;

	wire w74057;

	wire w78057;

	wire w82057;

	wire w86057;

	wire w90057;

	wire w169058;
	torch #(1'b0) c169058 (.i_clk(tick), .i_in(), .o_out(w169058));
	wire w173058;
	torch #(1'b0) c173058 (.i_clk(tick), .i_in(), .o_out(w173058));
	wire w177058;
	torch #(1'b0) c177058 (.i_clk(tick), .i_in(), .o_out(w177058));
	wire w181058;
	torch #(1'b0) c181058 (.i_clk(tick), .i_in(), .o_out(w181058));
	wire w185058;
	torch #(1'b0) c185058 (.i_clk(tick), .i_in(), .o_out(w185058));
	wire w189058;
	torch #(1'b0) c189058 (.i_clk(tick), .i_in(), .o_out(w189058));
	wire w193058;
	torch #(1'b0) c193058 (.i_clk(tick), .i_in(), .o_out(w193058));
	wire w170060;
	torch #(1'b1) c170060 (.i_clk(tick), .i_in(), .o_out(w170060));
	wire w174060;
	torch #(1'b1) c174060 (.i_clk(tick), .i_in(), .o_out(w174060));
	wire w178060;
	torch #(1'b1) c178060 (.i_clk(tick), .i_in(), .o_out(w178060));
	wire w182060;
	torch #(1'b1) c182060 (.i_clk(tick), .i_in(), .o_out(w182060));
	wire w186060;
	torch #(1'b1) c186060 (.i_clk(tick), .i_in(), .o_out(w186060));
	wire w190060;
	torch #(1'b1) c190060 (.i_clk(tick), .i_in(), .o_out(w190060));
	wire w194060;
	torch #(1'b1) c194060 (.i_clk(tick), .i_in(), .o_out(w194060));
	wire w47064;
	repeater #(1, 1'b1, 0, 0) c47064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47064));
	wire w81064;
	repeater #(1, 1'b1, 0, 0) c81064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81064));
	wire w172065;

	wire w197065;
	repeater #(2, 1'b0, 0, 0) c197065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197065));
	wire w192066;

	wire w47067;

	wire w81067;

	wire w48069;

	wire w82069;

	wire w176070;
	torch #(1'b1) c176070 (.i_clk(tick), .i_in(), .o_out(w176070));
	wire w180070;
	torch #(1'b1) c180070 (.i_clk(tick), .i_in(), .o_out(w180070));
	wire w184070;
	torch #(1'b1) c184070 (.i_clk(tick), .i_in(), .o_out(w184070));
	wire w188070;
	torch #(1'b1) c188070 (.i_clk(tick), .i_in(), .o_out(w188070));
	wire w47071;

	wire w48071;

	wire w81071;

	wire w82071;

	wire w169074;
	torch #(1'b0) c169074 (.i_clk(tick), .i_in(), .o_out(w169074));
	wire w173074;
	torch #(1'b0) c173074 (.i_clk(tick), .i_in(), .o_out(w173074));
	wire w177074;
	torch #(1'b0) c177074 (.i_clk(tick), .i_in(), .o_out(w177074));
	wire w181074;
	torch #(1'b0) c181074 (.i_clk(tick), .i_in(), .o_out(w181074));
	wire w185074;
	torch #(1'b0) c185074 (.i_clk(tick), .i_in(), .o_out(w185074));
	wire w189074;
	torch #(1'b0) c189074 (.i_clk(tick), .i_in(), .o_out(w189074));
	wire w193074;
	torch #(1'b0) c193074 (.i_clk(tick), .i_in(), .o_out(w193074));
	wire w105075;
	repeater #(1, 1'b1, 0, 0) c105075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105075));
	wire w157075;
	repeater #(1, 1'b1, 0, 0) c157075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157075));
	wire w111076;

	wire w115076;
	repeater #(1, 1'b1, 0, 0) c115076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115076));
	wire w147076;
	repeater #(1, 1'b1, 0, 0) c147076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147076));
	wire w151076;

	wire w170076;
	torch #(1'b1) c170076 (.i_clk(tick), .i_in(), .o_out(w170076));
	wire w174076;
	torch #(1'b1) c174076 (.i_clk(tick), .i_in(), .o_out(w174076));
	wire w178076;
	torch #(1'b1) c178076 (.i_clk(tick), .i_in(), .o_out(w178076));
	wire w182076;
	torch #(1'b1) c182076 (.i_clk(tick), .i_in(), .o_out(w182076));
	wire w186076;
	torch #(1'b1) c186076 (.i_clk(tick), .i_in(), .o_out(w186076));
	wire w190076;
	torch #(1'b1) c190076 (.i_clk(tick), .i_in(), .o_out(w190076));
	wire w194076;
	torch #(1'b1) c194076 (.i_clk(tick), .i_in(), .o_out(w194076));
	wire w56077;

	wire w57077;

	wire w90077;

	wire w91077;

	wire w112077;

	wire w150077;

	wire w111078;
	repeater #(2, 1'b0, 0, 0) c111078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111078));
	wire w151078;
	repeater #(2, 1'b1, 0, 0) c151078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151078));
	wire w105079;

	wire w106079;

	wire w156079;

	wire w157079;

	wire w104080;

	wire w113080;

	wire w149080;

	wire w158080;

	wire w172081;

	wire w197081;
	repeater #(2, 1'b0, 0, 0) c197081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197081));
	wire w192082;

	wire w37086;
	repeater #(1, 1'b0, 0, 0) c37086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37086));
	wire w45086;
	repeater #(1, 1'b0, 0, 0) c45086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45086));
	wire w53086;
	repeater #(1, 1'b0, 0, 0) c53086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53086));
	wire w71086;
	repeater #(1, 1'b0, 0, 0) c71086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71086));
	wire w79086;
	repeater #(1, 1'b0, 0, 0) c79086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79086));
	wire w87086;
	repeater #(1, 1'b0, 0, 0) c87086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87086));
	wire w176086;
	torch #(1'b1) c176086 (.i_clk(tick), .i_in(), .o_out(w176086));
	wire w180086;
	torch #(1'b1) c180086 (.i_clk(tick), .i_in(), .o_out(w180086));
	wire w184086;
	torch #(1'b1) c184086 (.i_clk(tick), .i_in(), .o_out(w184086));
	wire w188086;
	torch #(1'b1) c188086 (.i_clk(tick), .i_in(), .o_out(w188086));
	wire w37089;
	torch #(1'b0) c37089 (.i_clk(tick), .i_in(), .o_out(w37089));
	wire w45089;
	torch #(1'b0) c45089 (.i_clk(tick), .i_in(), .o_out(w45089));
	wire w53089;
	torch #(1'b0) c53089 (.i_clk(tick), .i_in(), .o_out(w53089));
	wire w71089;
	torch #(1'b0) c71089 (.i_clk(tick), .i_in(), .o_out(w71089));
	wire w79089;
	torch #(1'b0) c79089 (.i_clk(tick), .i_in(), .o_out(w79089));
	wire w87089;
	torch #(1'b0) c87089 (.i_clk(tick), .i_in(), .o_out(w87089));
	wire w33090;
	torch #(1'b0) c33090 (.i_clk(tick), .i_in(), .o_out(w33090));
	wire w41090;
	torch #(1'b0) c41090 (.i_clk(tick), .i_in(), .o_out(w41090));
	wire w49090;
	torch #(1'b0) c49090 (.i_clk(tick), .i_in(), .o_out(w49090));
	wire w57090;
	torch #(1'b0) c57090 (.i_clk(tick), .i_in(), .o_out(w57090));
	wire w67090;
	torch #(1'b0) c67090 (.i_clk(tick), .i_in(), .o_out(w67090));
	wire w75090;
	torch #(1'b0) c75090 (.i_clk(tick), .i_in(), .o_out(w75090));
	wire w83090;
	torch #(1'b0) c83090 (.i_clk(tick), .i_in(), .o_out(w83090));
	wire w91090;
	torch #(1'b0) c91090 (.i_clk(tick), .i_in(), .o_out(w91090));
	wire w169090;
	torch #(1'b0) c169090 (.i_clk(tick), .i_in(), .o_out(w169090));
	wire w173090;
	torch #(1'b0) c173090 (.i_clk(tick), .i_in(), .o_out(w173090));
	wire w177090;
	torch #(1'b0) c177090 (.i_clk(tick), .i_in(), .o_out(w177090));
	wire w181090;
	torch #(1'b0) c181090 (.i_clk(tick), .i_in(), .o_out(w181090));
	wire w185090;
	torch #(1'b0) c185090 (.i_clk(tick), .i_in(), .o_out(w185090));
	wire w189090;
	torch #(1'b0) c189090 (.i_clk(tick), .i_in(), .o_out(w189090));
	wire w193090;
	torch #(1'b0) c193090 (.i_clk(tick), .i_in(), .o_out(w193090));
	wire w170092;
	torch #(1'b1) c170092 (.i_clk(tick), .i_in(), .o_out(w170092));
	wire w174092;
	torch #(1'b1) c174092 (.i_clk(tick), .i_in(), .o_out(w174092));
	wire w178092;
	torch #(1'b1) c178092 (.i_clk(tick), .i_in(), .o_out(w178092));
	wire w182092;
	torch #(1'b1) c182092 (.i_clk(tick), .i_in(), .o_out(w182092));
	wire w186092;
	torch #(1'b1) c186092 (.i_clk(tick), .i_in(), .o_out(w186092));
	wire w190092;
	torch #(1'b1) c190092 (.i_clk(tick), .i_in(), .o_out(w190092));
	wire w194092;
	torch #(1'b1) c194092 (.i_clk(tick), .i_in(), .o_out(w194092));
	wire w172097;

	wire w197097;
	repeater #(2, 1'b0, 0, 0) c197097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197097));
	wire w192098;

	wire w1760102;
	torch #(1'b1) c1760102 (.i_clk(tick), .i_in(), .o_out(w1760102));
	wire w1800102;
	torch #(1'b1) c1800102 (.i_clk(tick), .i_in(), .o_out(w1800102));
	wire w1840102;
	torch #(1'b1) c1840102 (.i_clk(tick), .i_in(), .o_out(w1840102));
	wire w1880102;
	torch #(1'b1) c1880102 (.i_clk(tick), .i_in(), .o_out(w1880102));
	wire w1690106;
	torch #(1'b0) c1690106 (.i_clk(tick), .i_in(), .o_out(w1690106));
	wire w1730106;
	torch #(1'b0) c1730106 (.i_clk(tick), .i_in(), .o_out(w1730106));
	wire w1770106;
	torch #(1'b0) c1770106 (.i_clk(tick), .i_in(), .o_out(w1770106));
	wire w1810106;
	torch #(1'b0) c1810106 (.i_clk(tick), .i_in(), .o_out(w1810106));
	wire w1850106;
	torch #(1'b0) c1850106 (.i_clk(tick), .i_in(), .o_out(w1850106));
	wire w1890106;
	torch #(1'b0) c1890106 (.i_clk(tick), .i_in(), .o_out(w1890106));
	wire w1930106;
	torch #(1'b0) c1930106 (.i_clk(tick), .i_in(), .o_out(w1930106));
	wire w1700108;
	torch #(1'b1) c1700108 (.i_clk(tick), .i_in(), .o_out(w1700108));
	wire w1740108;
	torch #(1'b1) c1740108 (.i_clk(tick), .i_in(), .o_out(w1740108));
	wire w1780108;
	torch #(1'b1) c1780108 (.i_clk(tick), .i_in(), .o_out(w1780108));
	wire w1820108;
	torch #(1'b1) c1820108 (.i_clk(tick), .i_in(), .o_out(w1820108));
	wire w1860108;
	torch #(1'b1) c1860108 (.i_clk(tick), .i_in(), .o_out(w1860108));
	wire w1900108;
	torch #(1'b1) c1900108 (.i_clk(tick), .i_in(), .o_out(w1900108));
	wire w1940108;
	torch #(1'b1) c1940108 (.i_clk(tick), .i_in(), .o_out(w1940108));
	wire w1720113;

	wire w1970113;
	repeater #(2, 1'b0, 0, 0) c1970113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970113));
	wire w1920114;

	wire w1760118;
	torch #(1'b1) c1760118 (.i_clk(tick), .i_in(), .o_out(w1760118));
	wire w1800118;
	torch #(1'b1) c1800118 (.i_clk(tick), .i_in(), .o_out(w1800118));
	wire w1840118;
	torch #(1'b1) c1840118 (.i_clk(tick), .i_in(), .o_out(w1840118));
	wire w1880118;
	torch #(1'b1) c1880118 (.i_clk(tick), .i_in(), .o_out(w1880118));
	wire w1690122;
	torch #(1'b0) c1690122 (.i_clk(tick), .i_in(), .o_out(w1690122));
	wire w1730122;
	torch #(1'b0) c1730122 (.i_clk(tick), .i_in(), .o_out(w1730122));
	wire w1770122;
	torch #(1'b0) c1770122 (.i_clk(tick), .i_in(), .o_out(w1770122));
	wire w1810122;
	torch #(1'b0) c1810122 (.i_clk(tick), .i_in(), .o_out(w1810122));
	wire w1850122;
	torch #(1'b0) c1850122 (.i_clk(tick), .i_in(), .o_out(w1850122));
	wire w1890122;
	torch #(1'b0) c1890122 (.i_clk(tick), .i_in(), .o_out(w1890122));
	wire w1930122;
	torch #(1'b0) c1930122 (.i_clk(tick), .i_in(), .o_out(w1930122));
	wire w1700124;
	torch #(1'b1) c1700124 (.i_clk(tick), .i_in(), .o_out(w1700124));
	wire w1740124;
	torch #(1'b1) c1740124 (.i_clk(tick), .i_in(), .o_out(w1740124));
	wire w1780124;
	torch #(1'b1) c1780124 (.i_clk(tick), .i_in(), .o_out(w1780124));
	wire w1820124;
	torch #(1'b1) c1820124 (.i_clk(tick), .i_in(), .o_out(w1820124));
	wire w1860124;
	torch #(1'b1) c1860124 (.i_clk(tick), .i_in(), .o_out(w1860124));
	wire w1900124;
	torch #(1'b1) c1900124 (.i_clk(tick), .i_in(), .o_out(w1900124));
	wire w1940124;
	torch #(1'b1) c1940124 (.i_clk(tick), .i_in(), .o_out(w1940124));
	wire w1670136;
	repeater #(1, 1'b0, 0, 0) c1670136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1670136));
	wire w1710136;
	repeater #(1, 1'b0, 0, 0) c1710136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710136));
	wire w1750136;
	repeater #(1, 1'b0, 0, 0) c1750136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750136));
	wire w1790136;
	repeater #(1, 1'b0, 0, 0) c1790136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790136));
	wire w1830136;
	repeater #(1, 1'b0, 0, 0) c1830136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830136));
	wire w1870136;
	repeater #(1, 1'b0, 0, 0) c1870136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870136));
	wire w1910136;
	repeater #(1, 1'b0, 0, 0) c1910136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910136));
	wire w1680138;

	wire w1720138;

	wire w1760138;

	wire w1800138;

	wire w1840138;

	wire w1880138;

	wire w1920138;

	wire w1680139;

	wire w1720139;

	wire w1760139;

	wire w1800139;

	wire w1840139;

	wire w1880139;

	wire w1920139;

	wire w1670142;
	repeater #(1, 1'b1, 0, 0) c1670142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1670142));
	wire w1710142;
	repeater #(1, 1'b1, 0, 0) c1710142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710142));
	wire w1750142;
	repeater #(1, 1'b1, 0, 0) c1750142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750142));
	wire w1790142;
	repeater #(1, 1'b1, 0, 0) c1790142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790142));
	wire w1830142;
	repeater #(1, 1'b1, 0, 0) c1830142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830142));
	wire w1870142;
	repeater #(1, 1'b1, 0, 0) c1870142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1870142));
	wire w1910142;
	repeater #(1, 1'b1, 0, 0) c1910142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1910142));
	wire w1690143;

	wire w1730143;

	wire w1770143;

	wire w1810143;

	wire w1850143;

	wire w1890143;

	wire w1930143;

	wire w1680144;

	wire w1720144;

	wire w1760144;

	wire w1800144;

	wire w1840144;

	wire w1880144;

	wire w1920144;

	wire w1700146;
	torch #(1'b0) c1700146 (.i_clk(tick), .i_in(), .o_out(w1700146));
	wire w1740146;
	torch #(1'b0) c1740146 (.i_clk(tick), .i_in(), .o_out(w1740146));
	wire w1780146;
	torch #(1'b0) c1780146 (.i_clk(tick), .i_in(), .o_out(w1780146));
	wire w1820146;
	torch #(1'b0) c1820146 (.i_clk(tick), .i_in(), .o_out(w1820146));
	wire w1860146;
	torch #(1'b0) c1860146 (.i_clk(tick), .i_in(), .o_out(w1860146));
	wire w1900146;
	torch #(1'b0) c1900146 (.i_clk(tick), .i_in(), .o_out(w1900146));
	wire w1940146;
	torch #(1'b0) c1940146 (.i_clk(tick), .i_in(), .o_out(w1940146));
	wire w1700160;
	torch #(1'b0) c1700160 (.i_clk(tick), .i_in(), .o_out(w1700160));
	wire w1780160;
	torch #(1'b0) c1780160 (.i_clk(tick), .i_in(), .o_out(w1780160));
	wire w1860160;
	torch #(1'b0) c1860160 (.i_clk(tick), .i_in(), .o_out(w1860160));
	wire w1940160;
	torch #(1'b0) c1940160 (.i_clk(tick), .i_in(), .o_out(w1940160));
	wire w1700162;
	torch #(1'b0) c1700162 (.i_clk(tick), .i_in(), .o_out(w1700162));
	wire w1740162;
	torch #(1'b0) c1740162 (.i_clk(tick), .i_in(), .o_out(w1740162));
	wire w1860162;
	torch #(1'b0) c1860162 (.i_clk(tick), .i_in(), .o_out(w1860162));
	wire w1900162;
	torch #(1'b0) c1900162 (.i_clk(tick), .i_in(), .o_out(w1900162));
	wire w1700164;
	torch #(1'b0) c1700164 (.i_clk(tick), .i_in(), .o_out(w1700164));
	wire w1740164;
	torch #(1'b0) c1740164 (.i_clk(tick), .i_in(), .o_out(w1740164));
	wire w1780164;
	torch #(1'b0) c1780164 (.i_clk(tick), .i_in(), .o_out(w1780164));
	wire w1820164;
	torch #(1'b0) c1820164 (.i_clk(tick), .i_in(), .o_out(w1820164));
	wire w1700166;
	torch #(1'b0) c1700166 (.i_clk(tick), .i_in(), .o_out(w1700166));
	wire w1740166;
	torch #(1'b0) c1740166 (.i_clk(tick), .i_in(), .o_out(w1740166));
	wire w1780166;
	torch #(1'b0) c1780166 (.i_clk(tick), .i_in(), .o_out(w1780166));
	wire w1820166;
	torch #(1'b0) c1820166 (.i_clk(tick), .i_in(), .o_out(w1820166));
	wire w1860166;
	torch #(1'b0) c1860166 (.i_clk(tick), .i_in(), .o_out(w1860166));
	wire w1900166;
	torch #(1'b0) c1900166 (.i_clk(tick), .i_in(), .o_out(w1900166));
	wire w1940166;
	torch #(1'b0) c1940166 (.i_clk(tick), .i_in(), .o_out(w1940166));
	wire w1960166;
	torch #(1'b0) c1960166 (.i_clk(tick), .i_in(), .o_out(w1960166));
	wire w1980166;
	repeater #(1, 1'b0, 0, 0) c1980166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980166));
	wire w2000166;
	torch #(1'b0) c2000166 (.i_clk(tick), .i_in(), .o_out(w2000166));
	wire w5816;

	wire w9116;

	wire w9216;

	wire w12516;

	wire w12616;

	wire w15916;

	wire w16016;

	wire w19316;

	wire w5917;
	repeater #(1, 1'b1, 0, 0) c5917 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5917));
	wire w9317;
	repeater #(1, 1'b1, 0, 0) c9317 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9317));
	wire w12717;
	repeater #(1, 1'b1, 0, 0) c12717 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12717));
	wire w16117;
	repeater #(1, 1'b1, 0, 0) c16117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16117));
	wire w5618;

	wire w8918;

	wire w9018;

	wire w12318;

	wire w12418;

	wire w15718;

	wire w15818;

	wire w19118;

	wire w19418;
	repeater #(1, 1'b1, 0, 0) c19418 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19418));
	wire w5719;
	repeater #(1, 1'b1, 0, 0) c5719 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5719));
	wire w9119;
	repeater #(1, 1'b1, 0, 0) c9119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9119));
	wire w12519;
	repeater #(1, 1'b1, 0, 0) c12519 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w12519));
	wire w15919;
	repeater #(1, 1'b1, 0, 0) c15919 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15919));
	wire w19319;

	wire w54110;

	wire w87110;

	wire w88110;

	wire w121110;

	wire w122110;

	wire w155110;

	wire w156110;

	wire w189110;

	wire w192110;
	repeater #(1, 1'b1, 0, 0) c192110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192110));
	wire w55111;
	repeater #(1, 1'b1, 0, 0) c55111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55111));
	wire w89111;
	repeater #(1, 1'b1, 0, 0) c89111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89111));
	wire w123111;
	repeater #(1, 1'b1, 0, 0) c123111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123111));
	wire w157111;
	repeater #(1, 1'b1, 0, 0) c157111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157111));
	wire w191111;

	wire w52112;

	wire w85112;

	wire w86112;

	wire w119112;

	wire w120112;

	wire w153112;

	wire w154112;

	wire w187112;

	wire w190112;
	repeater #(1, 1'b1, 0, 0) c190112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190112));
	wire w53113;
	repeater #(1, 1'b1, 0, 0) c53113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w53113));
	wire w87113;
	repeater #(1, 1'b1, 0, 0) c87113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87113));
	wire w121113;
	repeater #(1, 1'b1, 0, 0) c121113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121113));
	wire w155113;
	repeater #(1, 1'b1, 0, 0) c155113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155113));
	wire w189113;

	wire w50114;

	wire w83114;

	wire w84114;

	wire w117114;

	wire w118114;

	wire w151114;

	wire w152114;

	wire w185114;

	wire w188114;
	repeater #(1, 1'b1, 0, 0) c188114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w188114));
	wire w51115;
	repeater #(1, 1'b1, 0, 0) c51115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51115));
	wire w85115;
	repeater #(1, 1'b1, 0, 0) c85115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85115));
	wire w119115;
	repeater #(1, 1'b1, 0, 0) c119115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119115));
	wire w153115;
	repeater #(1, 1'b1, 0, 0) c153115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153115));
	wire w187115;

	wire w48116;

	wire w81116;

	wire w82116;

	wire w115116;

	wire w116116;

	wire w149116;

	wire w150116;

	wire w183116;

	wire w186116;
	repeater #(1, 1'b1, 0, 0) c186116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186116));
	wire w49117;
	repeater #(1, 1'b1, 0, 0) c49117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49117));
	wire w83117;
	repeater #(1, 1'b1, 0, 0) c83117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83117));
	wire w117117;
	repeater #(1, 1'b1, 0, 0) c117117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117117));
	wire w151117;
	repeater #(1, 1'b1, 0, 0) c151117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151117));
	wire w185117;

	wire w46118;

	wire w79118;

	wire w80118;

	wire w113118;

	wire w114118;

	wire w147118;

	wire w148118;

	wire w181118;

	wire w184118;
	repeater #(1, 1'b1, 0, 0) c184118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184118));
	wire w47119;
	repeater #(1, 1'b1, 0, 0) c47119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47119));
	wire w81119;
	repeater #(1, 1'b1, 0, 0) c81119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81119));
	wire w115119;
	repeater #(1, 1'b1, 0, 0) c115119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115119));
	wire w149119;
	repeater #(1, 1'b1, 0, 0) c149119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149119));
	wire w183119;

	wire w44120;

	wire w77120;

	wire w78120;

	wire w111120;

	wire w112120;

	wire w145120;

	wire w146120;

	wire w179120;

	wire w182120;
	repeater #(1, 1'b1, 0, 0) c182120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182120));
	wire w45121;
	repeater #(1, 1'b1, 0, 0) c45121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45121));
	wire w79121;
	repeater #(1, 1'b1, 0, 0) c79121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79121));
	wire w113121;
	repeater #(1, 1'b1, 0, 0) c113121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113121));
	wire w147121;
	repeater #(1, 1'b1, 0, 0) c147121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147121));
	wire w181121;

	wire w42122;

	wire w75122;

	wire w76122;

	wire w109122;

	wire w110122;

	wire w143122;

	wire w144122;

	wire w177122;

	wire w180122;
	repeater #(1, 1'b1, 0, 0) c180122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180122));
	wire w43123;
	repeater #(1, 1'b1, 0, 0) c43123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w43123));
	wire w77123;
	repeater #(1, 1'b1, 0, 0) c77123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77123));
	wire w111123;
	repeater #(1, 1'b1, 0, 0) c111123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111123));
	wire w145123;
	repeater #(1, 1'b1, 0, 0) c145123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145123));
	wire w179123;

	wire w40124;

	wire w73124;

	wire w74124;

	wire w107124;

	wire w108124;

	wire w141124;

	wire w142124;

	wire w175124;

	wire w178124;
	repeater #(1, 1'b1, 0, 0) c178124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178124));
	wire w41125;
	repeater #(1, 1'b1, 0, 0) c41125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41125));
	wire w75125;
	repeater #(1, 1'b1, 0, 0) c75125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75125));
	wire w109125;
	repeater #(1, 1'b1, 0, 0) c109125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109125));
	wire w143125;
	repeater #(1, 1'b1, 0, 0) c143125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143125));
	wire w177125;

	wire w38126;

	wire w71126;

	wire w72126;

	wire w105126;

	wire w106126;

	wire w139126;

	wire w140126;

	wire w173126;

	wire w176126;
	repeater #(1, 1'b1, 0, 0) c176126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176126));
	wire w39127;
	repeater #(1, 1'b1, 0, 0) c39127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39127));
	wire w73127;
	repeater #(1, 1'b1, 0, 0) c73127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w73127));
	wire w107127;
	repeater #(1, 1'b1, 0, 0) c107127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107127));
	wire w141127;
	repeater #(1, 1'b1, 0, 0) c141127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141127));
	wire w175127;

	wire w36128;

	wire w69128;

	wire w70128;

	wire w103128;

	wire w104128;

	wire w137128;

	wire w138128;

	wire w171128;

	wire w174128;
	repeater #(1, 1'b1, 0, 0) c174128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174128));
	wire w37129;
	repeater #(1, 1'b1, 0, 0) c37129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37129));
	wire w71129;
	repeater #(1, 1'b1, 0, 0) c71129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71129));
	wire w105129;
	repeater #(1, 1'b1, 0, 0) c105129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105129));
	wire w139129;
	repeater #(1, 1'b1, 0, 0) c139129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139129));
	wire w173129;

	wire w34130;

	wire w67130;

	wire w68130;

	wire w101130;

	wire w102130;

	wire w135130;

	wire w136130;

	wire w169130;

	wire w172130;
	repeater #(1, 1'b1, 0, 0) c172130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172130));
	wire w35131;
	repeater #(1, 1'b1, 0, 0) c35131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35131));
	wire w69131;
	repeater #(1, 1'b1, 0, 0) c69131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69131));
	wire w103131;
	repeater #(1, 1'b1, 0, 0) c103131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103131));
	wire w137131;
	repeater #(1, 1'b1, 0, 0) c137131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137131));
	wire w171131;

	wire w65132;

	wire w99132;

	wire w133132;

	wire w167132;

	wire w170132;
	repeater #(1, 1'b1, 0, 0) c170132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170132));
	wire w33133;
	repeater #(1, 1'b1, 0, 0) c33133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33133));
	wire w67133;
	repeater #(1, 1'b1, 0, 0) c67133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67133));
	wire w101133;
	repeater #(1, 1'b1, 0, 0) c101133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101133));
	wire w135133;
	repeater #(1, 1'b1, 0, 0) c135133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135133));
	wire w169133;

	wire w168134;
	repeater #(2, 1'b1, 0, 0) c168134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168134));
	wire w170135;
	repeater #(1, 1'b1, 0, 0) c170135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170135));
	wire w169138;
	torch #(1'b1) c169138 (.i_clk(tick), .i_in(), .o_out(w169138));
	wire w173138;
	torch #(1'b1) c173138 (.i_clk(tick), .i_in(), .o_out(w173138));
	wire w177138;
	torch #(1'b1) c177138 (.i_clk(tick), .i_in(), .o_out(w177138));
	wire w181138;
	torch #(1'b1) c181138 (.i_clk(tick), .i_in(), .o_out(w181138));
	wire w185138;
	torch #(1'b1) c185138 (.i_clk(tick), .i_in(), .o_out(w185138));
	wire w189138;
	torch #(1'b1) c189138 (.i_clk(tick), .i_in(), .o_out(w189138));
	wire w193138;
	torch #(1'b1) c193138 (.i_clk(tick), .i_in(), .o_out(w193138));
	wire w38140;
	repeater #(1, 1'b1, 0, 0) c38140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38140));
	wire w72140;
	repeater #(1, 1'b1, 0, 0) c72140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72140));
	wire w170141;
	repeater #(1, 1'b1, 0, 0) c170141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170141));
	wire w174141;
	repeater #(1, 1'b1, 0, 0) c174141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174141));
	wire w178141;
	repeater #(1, 1'b1, 0, 0) c178141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178141));
	wire w182141;
	repeater #(1, 1'b1, 0, 0) c182141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182141));
	wire w186141;
	repeater #(1, 1'b1, 0, 0) c186141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186141));
	wire w190141;
	repeater #(1, 1'b1, 0, 0) c190141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190141));
	wire w194141;
	repeater #(1, 1'b1, 0, 0) c194141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194141));
	wire w169142;
	torch #(1'b1) c169142 (.i_clk(tick), .i_in(), .o_out(w169142));
	wire w173142;
	torch #(1'b1) c173142 (.i_clk(tick), .i_in(), .o_out(w173142));
	wire w177142;
	torch #(1'b1) c177142 (.i_clk(tick), .i_in(), .o_out(w177142));
	wire w181142;
	torch #(1'b1) c181142 (.i_clk(tick), .i_in(), .o_out(w181142));
	wire w185142;
	torch #(1'b1) c185142 (.i_clk(tick), .i_in(), .o_out(w185142));
	wire w189142;
	torch #(1'b1) c189142 (.i_clk(tick), .i_in(), .o_out(w189142));
	wire w193142;
	torch #(1'b1) c193142 (.i_clk(tick), .i_in(), .o_out(w193142));
	wire w38144;
	repeater #(1, 1'b1, 0, 0) c38144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38144));
	wire w72144;
	repeater #(1, 1'b1, 0, 0) c72144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72144));
	wire w168145;
	torch #(1'b0) c168145 (.i_clk(tick), .i_in(), .o_out(w168145));
	wire w172145;
	torch #(1'b0) c172145 (.i_clk(tick), .i_in(), .o_out(w172145));
	wire w176145;
	torch #(1'b0) c176145 (.i_clk(tick), .i_in(), .o_out(w176145));
	wire w180145;
	torch #(1'b0) c180145 (.i_clk(tick), .i_in(), .o_out(w180145));
	wire w184145;
	torch #(1'b0) c184145 (.i_clk(tick), .i_in(), .o_out(w184145));
	wire w188145;
	torch #(1'b0) c188145 (.i_clk(tick), .i_in(), .o_out(w188145));
	wire w192145;
	torch #(1'b0) c192145 (.i_clk(tick), .i_in(), .o_out(w192145));
	wire w101146;
	repeater #(1, 1'b1, 0, 0) c101146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101146));
	wire w105146;
	repeater #(1, 1'b1, 0, 0) c105146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105146));
	wire w109146;
	repeater #(1, 1'b1, 0, 0) c109146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109146));
	wire w113146;
	repeater #(1, 1'b0, 0, 0) c113146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113146));
	wire w117146;
	repeater #(1, 1'b1, 0, 0) c117146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w117146));
	wire w121146;
	repeater #(1, 1'b1, 0, 0) c121146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121146));
	wire w125146;
	repeater #(1, 1'b1, 0, 0) c125146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w125146));
	wire w137146;
	repeater #(1, 1'b1, 0, 0) c137146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137146));
	wire w141146;
	repeater #(1, 1'b1, 0, 0) c141146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w141146));
	wire w145146;
	repeater #(1, 1'b1, 0, 0) c145146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145146));
	wire w149146;
	repeater #(1, 1'b1, 0, 0) c149146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149146));
	wire w153146;
	repeater #(1, 1'b1, 0, 0) c153146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153146));
	wire w157146;
	repeater #(1, 1'b1, 0, 0) c157146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157146));
	wire w161146;
	repeater #(1, 1'b1, 0, 0) c161146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161146));
	wire w38147;

	wire w72147;

	wire w30149;

	wire w37149;

	wire w64149;

	wire w71149;

	wire w130156;
	repeater #(1, 1'b0, 0, 0) c130156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130156));
	wire w169160;
	torch #(1'b1) c169160 (.i_clk(tick), .i_in(), .o_out(w169160));
	wire w173160;
	torch #(1'b1) c173160 (.i_clk(tick), .i_in(), .o_out(w173160));
	wire w177160;
	torch #(1'b1) c177160 (.i_clk(tick), .i_in(), .o_out(w177160));
	wire w181160;
	torch #(1'b1) c181160 (.i_clk(tick), .i_in(), .o_out(w181160));
	wire w185160;
	torch #(1'b1) c185160 (.i_clk(tick), .i_in(), .o_out(w185160));
	wire w189160;
	torch #(1'b1) c189160 (.i_clk(tick), .i_in(), .o_out(w189160));
	wire w193160;
	torch #(1'b1) c193160 (.i_clk(tick), .i_in(), .o_out(w193160));
	wire w170161;
	repeater #(1, 1'b0, 0, 0) c170161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170161));
	wire w174161;
	repeater #(1, 1'b0, 0, 0) c174161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174161));
	wire w178161;
	repeater #(1, 1'b0, 0, 0) c178161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178161));
	wire w182161;
	repeater #(1, 1'b0, 0, 0) c182161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182161));
	wire w186161;
	repeater #(1, 1'b0, 0, 0) c186161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186161));
	wire w190161;
	repeater #(1, 1'b0, 0, 0) c190161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190161));
	wire w194161;
	repeater #(1, 1'b0, 0, 0) c194161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194161));
	wire w168163;

	wire w170163;
	repeater #(1, 1'b0, 0, 0) c170163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170163));
	wire w172163;

	wire w174163;
	repeater #(1, 1'b0, 0, 0) c174163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174163));
	wire w176163;

	wire w178163;
	repeater #(1, 1'b0, 0, 0) c178163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178163));
	wire w180163;

	wire w182163;
	repeater #(1, 1'b0, 0, 0) c182163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182163));
	wire w184163;

	wire w186163;
	repeater #(1, 1'b0, 0, 0) c186163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186163));
	wire w188163;

	wire w190163;
	repeater #(1, 1'b0, 0, 0) c190163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190163));
	wire w192163;

	wire w194163;
	repeater #(1, 1'b0, 0, 0) c194163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194163));
	wire w51164;
	repeater #(1, 1'b1, 0, 0) c51164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51164));
	wire w85164;
	repeater #(1, 1'b1, 0, 0) c85164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85164));
	wire w51167;

	wire w85167;

	wire w51171;

	wire w52171;

	wire w85171;

	wire w86171;

	wire w109175;

	wire w153175;

	wire w109176;
	repeater #(1, 1'b0, 0, 0) c109176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w109176));
	wire w153176;
	repeater #(1, 1'b1, 0, 0) c153176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153176));
	wire w169176;
	torch #(1'b1) c169176 (.i_clk(tick), .i_in(), .o_out(w169176));
	wire w173176;
	torch #(1'b1) c173176 (.i_clk(tick), .i_in(), .o_out(w173176));
	wire w177176;
	torch #(1'b1) c177176 (.i_clk(tick), .i_in(), .o_out(w177176));
	wire w181176;
	torch #(1'b1) c181176 (.i_clk(tick), .i_in(), .o_out(w181176));
	wire w185176;
	torch #(1'b1) c185176 (.i_clk(tick), .i_in(), .o_out(w185176));
	wire w189176;
	torch #(1'b1) c189176 (.i_clk(tick), .i_in(), .o_out(w189176));
	wire w193176;
	torch #(1'b1) c193176 (.i_clk(tick), .i_in(), .o_out(w193176));
	wire w170177;
	repeater #(1, 1'b0, 0, 0) c170177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170177));
	wire w174177;
	repeater #(1, 1'b0, 0, 0) c174177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174177));
	wire w178177;
	repeater #(1, 1'b0, 0, 0) c178177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178177));
	wire w182177;
	repeater #(1, 1'b0, 0, 0) c182177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182177));
	wire w186177;
	repeater #(1, 1'b0, 0, 0) c186177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186177));
	wire w190177;
	repeater #(1, 1'b0, 0, 0) c190177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190177));
	wire w194177;
	repeater #(1, 1'b0, 0, 0) c194177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194177));
	wire w110178;

	wire w114178;

	wire w148178;

	wire w152178;

	wire w110179;

	wire w112179;
	repeater #(1, 1'b0, 0, 0) c112179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112179));
	wire w113179;

	wire w149179;

	wire w150179;
	repeater #(1, 1'b1, 0, 0) c150179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150179));
	wire w152179;

	wire w168179;

	wire w170179;
	repeater #(1, 1'b0, 0, 0) c170179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170179));
	wire w172179;

	wire w174179;
	repeater #(1, 1'b0, 0, 0) c174179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174179));
	wire w176179;

	wire w178179;
	repeater #(1, 1'b0, 0, 0) c178179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178179));
	wire w180179;

	wire w182179;
	repeater #(1, 1'b0, 0, 0) c182179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182179));
	wire w184179;

	wire w186179;
	repeater #(1, 1'b0, 0, 0) c186179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186179));
	wire w188179;

	wire w190179;
	repeater #(1, 1'b0, 0, 0) c190179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190179));
	wire w192179;

	wire w194179;
	repeater #(1, 1'b0, 0, 0) c194179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194179));
	wire w47183;
	repeater #(2, 1'b0, 0, 0) c47183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47183));
	wire w50183;
	repeater #(2, 1'b0, 0, 0) c50183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50183));
	wire w54183;
	repeater #(1, 1'b0, 0, 0) c54183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54183));
	wire w69183;
	repeater #(1, 1'b0, 0, 0) c69183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69183));
	wire w74183;
	repeater #(2, 1'b0, 0, 0) c74183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74183));
	wire w76183;
	repeater #(2, 1'b0, 0, 0) c76183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76183));
	wire w78183;
	repeater #(2, 1'b0, 0, 0) c78183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78183));
	wire w45184;
	repeater #(1, 1'b0, 0, 0) c45184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w45184));
	wire w79184;
	repeater #(1, 1'b0, 0, 0) c79184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79184));
	wire w33186;
	repeater #(1, 1'b0, 0, 0) c33186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33186));
	wire w41186;
	repeater #(1, 1'b0, 0, 0) c41186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41186));
	wire w49186;
	repeater #(1, 1'b0, 0, 0) c49186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49186));
	wire w57186;
	repeater #(1, 1'b0, 0, 0) c57186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w57186));
	wire w67186;
	repeater #(1, 1'b0, 0, 0) c67186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w67186));
	wire w75186;
	repeater #(1, 1'b0, 0, 0) c75186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75186));
	wire w83186;
	repeater #(1, 1'b0, 0, 0) c83186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83186));
	wire w91186;
	repeater #(1, 1'b0, 0, 0) c91186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91186));
	wire w169192;
	torch #(1'b1) c169192 (.i_clk(tick), .i_in(), .o_out(w169192));
	wire w173192;
	torch #(1'b1) c173192 (.i_clk(tick), .i_in(), .o_out(w173192));
	wire w177192;
	torch #(1'b1) c177192 (.i_clk(tick), .i_in(), .o_out(w177192));
	wire w181192;
	torch #(1'b1) c181192 (.i_clk(tick), .i_in(), .o_out(w181192));
	wire w185192;
	torch #(1'b1) c185192 (.i_clk(tick), .i_in(), .o_out(w185192));
	wire w189192;
	torch #(1'b1) c189192 (.i_clk(tick), .i_in(), .o_out(w189192));
	wire w193192;
	torch #(1'b1) c193192 (.i_clk(tick), .i_in(), .o_out(w193192));
	wire w170193;
	repeater #(1, 1'b0, 0, 0) c170193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170193));
	wire w174193;
	repeater #(1, 1'b0, 0, 0) c174193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174193));
	wire w178193;
	repeater #(1, 1'b0, 0, 0) c178193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178193));
	wire w182193;
	repeater #(1, 1'b0, 0, 0) c182193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182193));
	wire w186193;
	repeater #(1, 1'b0, 0, 0) c186193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186193));
	wire w190193;
	repeater #(1, 1'b0, 0, 0) c190193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190193));
	wire w194193;
	repeater #(1, 1'b0, 0, 0) c194193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194193));
	wire w47194;

	wire w81194;

	wire w39195;

	wire w43195;

	wire w46195;

	wire w48195;

	wire w51195;

	wire w73195;

	wire w77195;

	wire w80195;

	wire w82195;

	wire w85195;

	wire w168195;

	wire w170195;
	repeater #(1, 1'b0, 0, 0) c170195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170195));
	wire w172195;

	wire w174195;
	repeater #(1, 1'b0, 0, 0) c174195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174195));
	wire w176195;

	wire w178195;
	repeater #(1, 1'b0, 0, 0) c178195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178195));
	wire w180195;

	wire w182195;
	repeater #(1, 1'b0, 0, 0) c182195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182195));
	wire w184195;

	wire w186195;
	repeater #(1, 1'b0, 0, 0) c186195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186195));
	wire w188195;

	wire w190195;
	repeater #(1, 1'b0, 0, 0) c190195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190195));
	wire w192195;

	wire w194195;
	repeater #(1, 1'b0, 0, 0) c194195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194195));
	wire w38196;

	wire w40196;

	wire w42196;

	wire w44196;

	wire w47196;

	wire w50196;

	wire w52196;

	wire w72196;

	wire w74196;

	wire w76196;

	wire w78196;

	wire w81196;

	wire w84196;

	wire w86196;

	wire w43197;

	wire w77197;

	wire w39198;

	wire w43198;

	wire w44198;

	wire w48198;

	wire w50198;

	wire w52198;

	wire w73198;

	wire w77198;

	wire w78198;

	wire w82198;

	wire w84198;

	wire w86198;

	wire w1731108;
	torch #(1'b1) c1731108 (.i_clk(tick), .i_in(), .o_out(w1731108));
	wire w1771108;
	torch #(1'b1) c1771108 (.i_clk(tick), .i_in(), .o_out(w1771108));
	wire w1811108;
	torch #(1'b1) c1811108 (.i_clk(tick), .i_in(), .o_out(w1811108));
	wire w1851108;
	torch #(1'b1) c1851108 (.i_clk(tick), .i_in(), .o_out(w1851108));
	wire w1891108;
	torch #(1'b1) c1891108 (.i_clk(tick), .i_in(), .o_out(w1891108));
	wire w1931108;
	torch #(1'b1) c1931108 (.i_clk(tick), .i_in(), .o_out(w1931108));
	wire w1701109;
	repeater #(1, 1'b0, 0, 0) c1701109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701109));
	wire w1741109;
	repeater #(1, 1'b0, 0, 0) c1741109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741109));
	wire w1781109;
	repeater #(1, 1'b0, 0, 0) c1781109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781109));
	wire w1821109;
	repeater #(1, 1'b0, 0, 0) c1821109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821109));
	wire w1861109;
	repeater #(1, 1'b0, 0, 0) c1861109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861109));
	wire w1901109;
	repeater #(1, 1'b0, 0, 0) c1901109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901109));
	wire w1941109;
	repeater #(1, 1'b0, 0, 0) c1941109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941109));
	wire w1681111;

	wire w1701111;
	repeater #(1, 1'b0, 0, 0) c1701111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701111));
	wire w1721111;

	wire w1741111;
	repeater #(1, 1'b0, 0, 0) c1741111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741111));
	wire w1761111;

	wire w1781111;
	repeater #(1, 1'b0, 0, 0) c1781111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781111));
	wire w1801111;

	wire w1821111;
	repeater #(1, 1'b0, 0, 0) c1821111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821111));
	wire w1841111;

	wire w1861111;
	repeater #(1, 1'b0, 0, 0) c1861111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861111));
	wire w1881111;

	wire w1901111;
	repeater #(1, 1'b0, 0, 0) c1901111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901111));
	wire w1921111;

	wire w1941111;
	repeater #(1, 1'b0, 0, 0) c1941111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941111));
	wire w1691124;
	torch #(1'b1) c1691124 (.i_clk(tick), .i_in(), .o_out(w1691124));
	wire w1731124;
	torch #(1'b1) c1731124 (.i_clk(tick), .i_in(), .o_out(w1731124));
	wire w1771124;
	torch #(1'b1) c1771124 (.i_clk(tick), .i_in(), .o_out(w1771124));
	wire w1811124;
	torch #(1'b1) c1811124 (.i_clk(tick), .i_in(), .o_out(w1811124));
	wire w1851124;
	torch #(1'b1) c1851124 (.i_clk(tick), .i_in(), .o_out(w1851124));
	wire w1891124;
	torch #(1'b1) c1891124 (.i_clk(tick), .i_in(), .o_out(w1891124));
	wire w1931124;
	torch #(1'b1) c1931124 (.i_clk(tick), .i_in(), .o_out(w1931124));
	wire w1701125;
	repeater #(1, 1'b0, 0, 0) c1701125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701125));
	wire w1741125;
	repeater #(1, 1'b0, 0, 0) c1741125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741125));
	wire w1781125;
	repeater #(1, 1'b0, 0, 0) c1781125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781125));
	wire w1821125;
	repeater #(1, 1'b0, 0, 0) c1821125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821125));
	wire w1861125;
	repeater #(1, 1'b0, 0, 0) c1861125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861125));
	wire w1901125;
	repeater #(1, 1'b0, 0, 0) c1901125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901125));
	wire w1941125;
	repeater #(1, 1'b0, 0, 0) c1941125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941125));
	wire w1681127;

	wire w1701127;
	repeater #(1, 1'b0, 0, 0) c1701127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701127));
	wire w1721127;

	wire w1741127;
	repeater #(1, 1'b0, 0, 0) c1741127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741127));
	wire w1761127;

	wire w1781127;
	repeater #(1, 1'b0, 0, 0) c1781127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781127));
	wire w1801127;

	wire w1821127;
	repeater #(1, 1'b0, 0, 0) c1821127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821127));
	wire w1841127;

	wire w1861127;
	repeater #(1, 1'b0, 0, 0) c1861127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861127));
	wire w1881127;

	wire w1901127;
	repeater #(1, 1'b0, 0, 0) c1901127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901127));
	wire w1921127;

	wire w1941127;
	repeater #(1, 1'b0, 0, 0) c1941127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941127));
	wire w1691133;
	torch #(1'b1) c1691133 (.i_clk(tick), .i_in(), .o_out(w1691133));
	wire w1731133;
	torch #(1'b1) c1731133 (.i_clk(tick), .i_in(), .o_out(w1731133));
	wire w1771133;
	torch #(1'b1) c1771133 (.i_clk(tick), .i_in(), .o_out(w1771133));
	wire w1811133;
	torch #(1'b1) c1811133 (.i_clk(tick), .i_in(), .o_out(w1811133));
	wire w1851133;
	torch #(1'b1) c1851133 (.i_clk(tick), .i_in(), .o_out(w1851133));
	wire w1891133;
	torch #(1'b1) c1891133 (.i_clk(tick), .i_in(), .o_out(w1891133));
	wire w1931133;
	torch #(1'b1) c1931133 (.i_clk(tick), .i_in(), .o_out(w1931133));
	wire w15409;
	repeater #(1, 1'b0, 0, 0) c15409 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15409));
	wire w15809;
	repeater #(1, 1'b0, 0, 0) c15809 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15809));
	wire w16209;
	repeater #(1, 1'b0, 0, 0) c16209 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16209));
	wire w16609;
	repeater #(1, 1'b0, 0, 0) c16609 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16609));
	wire w17009;
	repeater #(1, 1'b0, 0, 0) c17009 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17009));
	wire w17409;
	repeater #(1, 1'b0, 0, 0) c17409 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17409));
	wire w17809;
	repeater #(1, 1'b0, 0, 0) c17809 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17809));
	wire w153010;
	repeater #(1, 1'b1, 0, 0) c153010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153010));
	wire w157010;
	repeater #(1, 1'b1, 0, 0) c157010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w157010));
	wire w161010;
	repeater #(1, 1'b1, 0, 0) c161010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161010));
	wire w165010;
	repeater #(1, 1'b1, 0, 0) c165010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w165010));
	wire w169010;
	repeater #(1, 1'b1, 0, 0) c169010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169010));
	wire w173010;
	repeater #(1, 1'b1, 0, 0) c173010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w173010));
	wire w177010;
	repeater #(1, 1'b1, 0, 0) c177010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177010));
	wire w154019;
	repeater #(1, 1'b0, 0, 0) c154019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154019));
	wire w158019;
	repeater #(1, 1'b0, 0, 0) c158019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158019));
	wire w162019;
	repeater #(1, 1'b0, 0, 0) c162019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162019));
	wire w166019;
	repeater #(1, 1'b0, 0, 0) c166019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166019));
	wire w170019;
	repeater #(1, 1'b0, 0, 0) c170019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170019));
	wire w174019;
	repeater #(1, 1'b0, 0, 0) c174019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174019));
	wire w178019;
	repeater #(1, 1'b0, 0, 0) c178019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178019));
	wire w164023;
	repeater #(1, 1'b0, 0, 0) c164023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164023));
	wire w182023;
	repeater #(2, 1'b0, 0, 0) c182023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182023));
	wire w164025;
	repeater #(1, 1'b0, 0, 0) c164025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164025));
	wire w182025;
	repeater #(2, 1'b0, 0, 0) c182025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182025));
	wire w164027;
	repeater #(1, 1'b0, 0, 0) c164027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164027));
	wire w182027;
	repeater #(1, 1'b0, 0, 0) c182027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182027));
	wire w164029;
	repeater #(1, 1'b0, 0, 0) c164029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164029));
	wire w182029;
	repeater #(2, 1'b0, 0, 0) c182029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182029));
	wire w153044;
	torch #(1'b1) c153044 (.i_clk(tick), .i_in(), .o_out(w153044));
	wire w157044;
	torch #(1'b1) c157044 (.i_clk(tick), .i_in(), .o_out(w157044));
	wire w161044;
	torch #(1'b1) c161044 (.i_clk(tick), .i_in(), .o_out(w161044));
	wire w165044;
	torch #(1'b1) c165044 (.i_clk(tick), .i_in(), .o_out(w165044));
	wire w169044;
	torch #(1'b1) c169044 (.i_clk(tick), .i_in(), .o_out(w169044));
	wire w173044;
	torch #(1'b1) c173044 (.i_clk(tick), .i_in(), .o_out(w173044));
	wire w177044;
	torch #(1'b1) c177044 (.i_clk(tick), .i_in(), .o_out(w177044));
	wire w61049;

	wire w95049;

	wire w129049;

	wire w163049;

	wire w60050;
	repeater #(1, 1'b1, 0, 0) c60050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60050));
	wire w94050;
	repeater #(1, 1'b1, 0, 0) c94050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94050));
	wire w128050;
	repeater #(1, 1'b1, 0, 0) c128050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128050));
	wire w162050;
	repeater #(1, 1'b1, 0, 0) c162050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162050));
	wire w59051;

	wire w93051;

	wire w127051;

	wire w161051;

	wire w58052;
	repeater #(1, 1'b1, 0, 0) c58052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58052));
	wire w92052;
	repeater #(1, 1'b1, 0, 0) c92052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92052));
	wire w126052;
	repeater #(1, 1'b1, 0, 0) c126052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126052));
	wire w160052;
	repeater #(1, 1'b1, 0, 0) c160052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160052));
	wire w57053;

	wire w91053;

	wire w125053;

	wire w159053;

	wire w56054;
	repeater #(1, 1'b1, 0, 0) c56054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56054));
	wire w90054;
	repeater #(1, 1'b1, 0, 0) c90054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90054));
	wire w124054;
	repeater #(1, 1'b1, 0, 0) c124054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124054));
	wire w158054;
	repeater #(1, 1'b1, 0, 0) c158054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158054));
	wire w55055;

	wire w89055;

	wire w123055;

	wire w157055;

	wire w54056;
	repeater #(1, 1'b1, 0, 0) c54056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54056));
	wire w88056;
	repeater #(1, 1'b1, 0, 0) c88056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88056));
	wire w122056;
	repeater #(1, 1'b1, 0, 0) c122056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122056));
	wire w156056;
	repeater #(1, 1'b1, 0, 0) c156056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156056));
	wire w53057;

	wire w87057;

	wire w121057;

	wire w155057;

	wire w52058;
	repeater #(1, 1'b1, 0, 0) c52058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52058));
	wire w86058;
	repeater #(1, 1'b1, 0, 0) c86058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86058));
	wire w120058;
	repeater #(1, 1'b1, 0, 0) c120058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120058));
	wire w154058;
	repeater #(1, 1'b1, 0, 0) c154058 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154058));
	wire w51059;

	wire w85059;

	wire w119059;

	wire w153059;

	wire w50060;
	repeater #(1, 1'b1, 0, 0) c50060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50060));
	wire w84060;
	repeater #(1, 1'b1, 0, 0) c84060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84060));
	wire w118060;
	repeater #(1, 1'b1, 0, 0) c118060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w118060));
	wire w152060;
	repeater #(1, 1'b1, 0, 0) c152060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152060));
	wire w49061;

	wire w83061;

	wire w117061;

	wire w151061;

	wire w48062;
	repeater #(1, 1'b1, 0, 0) c48062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48062));
	wire w82062;
	repeater #(1, 1'b1, 0, 0) c82062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82062));
	wire w116062;
	repeater #(1, 1'b1, 0, 0) c116062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116062));
	wire w150062;
	repeater #(1, 1'b1, 0, 0) c150062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150062));
	wire w47063;

	wire w81063;

	wire w115063;

	wire w149063;

	wire w46064;
	repeater #(1, 1'b1, 0, 0) c46064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46064));
	wire w80064;
	repeater #(1, 1'b1, 0, 0) c80064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80064));
	wire w114064;
	repeater #(1, 1'b1, 0, 0) c114064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114064));
	wire w148064;
	repeater #(1, 1'b1, 0, 0) c148064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148064));
	wire w45065;

	wire w79065;

	wire w113065;

	wire w147065;

	wire w44066;
	repeater #(1, 1'b1, 0, 0) c44066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w44066));
	wire w78066;
	repeater #(1, 1'b1, 0, 0) c78066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78066));
	wire w112066;
	repeater #(1, 1'b1, 0, 0) c112066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112066));
	wire w146066;
	repeater #(1, 1'b1, 0, 0) c146066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146066));
	wire w43067;

	wire w77067;

	wire w111067;

	wire w145067;

	wire w42068;
	repeater #(1, 1'b1, 0, 0) c42068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42068));
	wire w76068;
	repeater #(1, 1'b1, 0, 0) c76068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76068));
	wire w110068;
	repeater #(1, 1'b1, 0, 0) c110068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110068));
	wire w144068;
	repeater #(1, 1'b1, 0, 0) c144068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144068));
	wire w41069;

	wire w75069;

	wire w109069;

	wire w143069;

	wire w40070;
	repeater #(1, 1'b1, 0, 0) c40070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40070));
	wire w74070;
	repeater #(1, 1'b1, 0, 0) c74070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74070));
	wire w108070;
	repeater #(1, 1'b1, 0, 0) c108070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108070));
	wire w142070;
	repeater #(1, 1'b1, 0, 0) c142070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142070));
	wire w39071;

	wire w73071;

	wire w107071;

	wire w141071;

	wire w38072;
	repeater #(1, 1'b1, 0, 0) c38072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38072));
	wire w72072;
	repeater #(1, 1'b1, 0, 0) c72072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72072));
	wire w106072;
	repeater #(1, 1'b1, 0, 0) c106072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106072));
	wire w140072;
	repeater #(1, 1'b1, 0, 0) c140072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140072));
	wire w37073;

	wire w71073;

	wire w105073;

	wire w139073;

	wire w36074;
	repeater #(1, 1'b1, 0, 0) c36074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36074));
	wire w70074;
	repeater #(1, 1'b1, 0, 0) c70074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70074));
	wire w104074;
	repeater #(1, 1'b1, 0, 0) c104074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104074));
	wire w138074;
	repeater #(1, 1'b1, 0, 0) c138074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138074));
	wire w35075;

	wire w69075;

	wire w103075;

	wire w137075;

	wire w34076;
	repeater #(1, 1'b1, 0, 0) c34076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34076));
	wire w68076;
	repeater #(1, 1'b1, 0, 0) c68076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68076));
	wire w102076;
	repeater #(1, 1'b1, 0, 0) c102076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102076));
	wire w136076;
	repeater #(1, 1'b1, 0, 0) c136076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136076));
	wire w85080;
	torch #(1'b0) c85080 (.i_clk(tick), .i_in(), .o_out(w85080));
	wire w89080;
	torch #(1'b0) c89080 (.i_clk(tick), .i_in(), .o_out(w89080));
	wire w93080;
	torch #(1'b0) c93080 (.i_clk(tick), .i_in(), .o_out(w93080));
	wire w97080;
	torch #(1'b1) c97080 (.i_clk(tick), .i_in(), .o_out(w97080));
	wire w101080;
	torch #(1'b0) c101080 (.i_clk(tick), .i_in(), .o_out(w101080));
	wire w105080;
	torch #(1'b0) c105080 (.i_clk(tick), .i_in(), .o_out(w105080));
	wire w109080;
	torch #(1'b0) c109080 (.i_clk(tick), .i_in(), .o_out(w109080));
	wire w121080;
	torch #(1'b0) c121080 (.i_clk(tick), .i_in(), .o_out(w121080));
	wire w125080;
	torch #(1'b0) c125080 (.i_clk(tick), .i_in(), .o_out(w125080));
	wire w129080;
	torch #(1'b0) c129080 (.i_clk(tick), .i_in(), .o_out(w129080));
	wire w133080;
	torch #(1'b0) c133080 (.i_clk(tick), .i_in(), .o_out(w133080));
	wire w137080;
	torch #(1'b0) c137080 (.i_clk(tick), .i_in(), .o_out(w137080));
	wire w141080;
	torch #(1'b0) c141080 (.i_clk(tick), .i_in(), .o_out(w141080));
	wire w145080;
	torch #(1'b0) c145080 (.i_clk(tick), .i_in(), .o_out(w145080));
	wire w152082;
	repeater #(1, 1'b1, 0, 0) c152082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152082));
	wire w156082;
	repeater #(1, 1'b1, 0, 0) c156082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156082));
	wire w160082;
	repeater #(1, 1'b1, 0, 0) c160082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160082));
	wire w164082;
	repeater #(1, 1'b1, 0, 0) c164082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164082));
	wire w168082;
	repeater #(1, 1'b1, 0, 0) c168082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168082));
	wire w172082;
	repeater #(1, 1'b1, 0, 0) c172082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172082));
	wire w176082;
	repeater #(1, 1'b1, 0, 0) c176082 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176082));
	wire w18083;
	repeater #(1, 1'b1, 0, 0) c18083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18083));
	wire w52083;
	repeater #(1, 1'b1, 0, 0) c52083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52083));
	wire w152083;
	repeater #(1, 1'b1, 0, 0) c152083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152083));
	wire w154083;
	repeater #(1, 1'b0, 0, 0) c154083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154083));
	wire w156083;
	repeater #(1, 1'b1, 0, 0) c156083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w156083));
	wire w158083;
	repeater #(1, 1'b0, 0, 0) c158083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158083));
	wire w160083;
	repeater #(1, 1'b1, 0, 0) c160083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160083));
	wire w162083;
	repeater #(1, 1'b0, 0, 0) c162083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162083));
	wire w164083;
	repeater #(1, 1'b1, 0, 0) c164083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164083));
	wire w166083;
	repeater #(1, 1'b0, 0, 0) c166083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166083));
	wire w168083;
	repeater #(1, 1'b1, 0, 0) c168083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168083));
	wire w170083;
	repeater #(1, 1'b0, 0, 0) c170083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170083));
	wire w172083;
	repeater #(1, 1'b1, 0, 0) c172083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172083));
	wire w174083;
	repeater #(1, 1'b0, 0, 0) c174083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174083));
	wire w176083;
	repeater #(1, 1'b1, 0, 0) c176083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176083));
	wire w178083;
	repeater #(1, 1'b0, 0, 0) c178083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178083));
	wire w153084;
	torch #(1'b0) c153084 (.i_clk(tick), .i_in(), .o_out(w153084));
	wire w157084;
	torch #(1'b0) c157084 (.i_clk(tick), .i_in(), .o_out(w157084));
	wire w161084;
	torch #(1'b0) c161084 (.i_clk(tick), .i_in(), .o_out(w161084));
	wire w165084;
	torch #(1'b0) c165084 (.i_clk(tick), .i_in(), .o_out(w165084));
	wire w169084;
	torch #(1'b0) c169084 (.i_clk(tick), .i_in(), .o_out(w169084));
	wire w173084;
	torch #(1'b0) c173084 (.i_clk(tick), .i_in(), .o_out(w173084));
	wire w177084;
	torch #(1'b0) c177084 (.i_clk(tick), .i_in(), .o_out(w177084));
	wire w18087;
	repeater #(1, 1'b1, 0, 0) c18087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18087));
	wire w52087;
	repeater #(1, 1'b1, 0, 0) c52087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52087));
	wire w18090;

	wire w52090;

	wire w147092;
	repeater #(2, 1'b0, 0, 0) c147092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147092));
	wire w17093;

	wire w51093;

	wire w154094;

	wire w158094;

	wire w162094;

	wire w166094;

	wire w170094;

	wire w174094;

	wire w178094;

	wire w113098;

	wire w1550103;
	torch #(1'b1) c1550103 (.i_clk(tick), .i_in(), .o_out(w1550103));
	wire w1590103;
	torch #(1'b1) c1590103 (.i_clk(tick), .i_in(), .o_out(w1590103));
	wire w1630103;
	torch #(1'b1) c1630103 (.i_clk(tick), .i_in(), .o_out(w1630103));
	wire w1670103;
	torch #(1'b1) c1670103 (.i_clk(tick), .i_in(), .o_out(w1670103));
	wire w1710103;
	torch #(1'b1) c1710103 (.i_clk(tick), .i_in(), .o_out(w1710103));
	wire w1750103;
	torch #(1'b1) c1750103 (.i_clk(tick), .i_in(), .o_out(w1750103));
	wire w1790103;
	torch #(1'b1) c1790103 (.i_clk(tick), .i_in(), .o_out(w1790103));
	wire w1470105;
	repeater #(1, 1'b0, 0, 0) c1470105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470105));
	wire w1540105;
	torch #(1'b0) c1540105 (.i_clk(tick), .i_in(), .o_out(w1540105));
	wire w1580105;
	torch #(1'b0) c1580105 (.i_clk(tick), .i_in(), .o_out(w1580105));
	wire w1620105;
	torch #(1'b0) c1620105 (.i_clk(tick), .i_in(), .o_out(w1620105));
	wire w1660105;
	torch #(1'b0) c1660105 (.i_clk(tick), .i_in(), .o_out(w1660105));
	wire w1700105;
	torch #(1'b0) c1700105 (.i_clk(tick), .i_in(), .o_out(w1700105));
	wire w1740105;
	torch #(1'b0) c1740105 (.i_clk(tick), .i_in(), .o_out(w1740105));
	wire w1780105;
	torch #(1'b0) c1780105 (.i_clk(tick), .i_in(), .o_out(w1780105));
	wire w1470106;
	repeater #(1, 1'b0, 0, 0) c1470106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470106));
	wire w1470107;
	repeater #(1, 1'b0, 0, 0) c1470107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470107));
	wire w1540110;

	wire w1580110;

	wire w1620110;

	wire w1660110;

	wire w1700110;

	wire w1740110;

	wire w1780110;

	wire w1550119;
	torch #(1'b1) c1550119 (.i_clk(tick), .i_in(), .o_out(w1550119));
	wire w1590119;
	torch #(1'b1) c1590119 (.i_clk(tick), .i_in(), .o_out(w1590119));
	wire w1630119;
	torch #(1'b1) c1630119 (.i_clk(tick), .i_in(), .o_out(w1630119));
	wire w1670119;
	torch #(1'b1) c1670119 (.i_clk(tick), .i_in(), .o_out(w1670119));
	wire w1710119;
	torch #(1'b1) c1710119 (.i_clk(tick), .i_in(), .o_out(w1710119));
	wire w1750119;
	torch #(1'b1) c1750119 (.i_clk(tick), .i_in(), .o_out(w1750119));
	wire w1790119;
	torch #(1'b1) c1790119 (.i_clk(tick), .i_in(), .o_out(w1790119));
	wire w1470121;
	repeater #(1, 1'b0, 0, 0) c1470121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470121));
	wire w1540121;
	torch #(1'b0) c1540121 (.i_clk(tick), .i_in(), .o_out(w1540121));
	wire w1580121;
	torch #(1'b0) c1580121 (.i_clk(tick), .i_in(), .o_out(w1580121));
	wire w1620121;
	torch #(1'b0) c1620121 (.i_clk(tick), .i_in(), .o_out(w1620121));
	wire w1660121;
	torch #(1'b0) c1660121 (.i_clk(tick), .i_in(), .o_out(w1660121));
	wire w1700121;
	torch #(1'b0) c1700121 (.i_clk(tick), .i_in(), .o_out(w1700121));
	wire w1740121;
	torch #(1'b0) c1740121 (.i_clk(tick), .i_in(), .o_out(w1740121));
	wire w1780121;
	torch #(1'b0) c1780121 (.i_clk(tick), .i_in(), .o_out(w1780121));
	wire w1470122;
	repeater #(1, 1'b0, 0, 0) c1470122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470122));
	wire w1470123;
	repeater #(1, 1'b0, 0, 0) c1470123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470123));
	wire w1540126;

	wire w1580126;

	wire w1620126;

	wire w1660126;

	wire w1700126;

	wire w1740126;

	wire w1780126;

	wire w1550135;
	torch #(1'b1) c1550135 (.i_clk(tick), .i_in(), .o_out(w1550135));
	wire w1590135;
	torch #(1'b1) c1590135 (.i_clk(tick), .i_in(), .o_out(w1590135));
	wire w1630135;
	torch #(1'b1) c1630135 (.i_clk(tick), .i_in(), .o_out(w1630135));
	wire w1670135;
	torch #(1'b1) c1670135 (.i_clk(tick), .i_in(), .o_out(w1670135));
	wire w1710135;
	torch #(1'b1) c1710135 (.i_clk(tick), .i_in(), .o_out(w1710135));
	wire w1750135;
	torch #(1'b1) c1750135 (.i_clk(tick), .i_in(), .o_out(w1750135));
	wire w1790135;
	torch #(1'b1) c1790135 (.i_clk(tick), .i_in(), .o_out(w1790135));
	wire w1470137;
	repeater #(1, 1'b0, 0, 0) c1470137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470137));
	wire w1540137;
	torch #(1'b0) c1540137 (.i_clk(tick), .i_in(), .o_out(w1540137));
	wire w1580137;
	torch #(1'b0) c1580137 (.i_clk(tick), .i_in(), .o_out(w1580137));
	wire w1620137;
	torch #(1'b0) c1620137 (.i_clk(tick), .i_in(), .o_out(w1620137));
	wire w1660137;
	torch #(1'b0) c1660137 (.i_clk(tick), .i_in(), .o_out(w1660137));
	wire w1700137;
	torch #(1'b0) c1700137 (.i_clk(tick), .i_in(), .o_out(w1700137));
	wire w1740137;
	torch #(1'b0) c1740137 (.i_clk(tick), .i_in(), .o_out(w1740137));
	wire w1780137;
	torch #(1'b0) c1780137 (.i_clk(tick), .i_in(), .o_out(w1780137));
	wire w1470138;
	repeater #(1, 1'b0, 0, 0) c1470138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470138));
	wire w1470139;
	repeater #(1, 1'b0, 0, 0) c1470139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470139));
	wire w1540142;

	wire w1580142;

	wire w1620142;

	wire w1660142;

	wire w1700142;

	wire w1740142;

	wire w1780142;

	wire w1550151;
	torch #(1'b1) c1550151 (.i_clk(tick), .i_in(), .o_out(w1550151));
	wire w1590151;
	torch #(1'b1) c1590151 (.i_clk(tick), .i_in(), .o_out(w1590151));
	wire w1630151;
	torch #(1'b1) c1630151 (.i_clk(tick), .i_in(), .o_out(w1630151));
	wire w1670151;
	torch #(1'b1) c1670151 (.i_clk(tick), .i_in(), .o_out(w1670151));
	wire w1710151;
	torch #(1'b1) c1710151 (.i_clk(tick), .i_in(), .o_out(w1710151));
	wire w1750151;
	torch #(1'b1) c1750151 (.i_clk(tick), .i_in(), .o_out(w1750151));
	wire w1790151;
	torch #(1'b1) c1790151 (.i_clk(tick), .i_in(), .o_out(w1790151));
	wire w1470153;
	repeater #(1, 1'b0, 0, 0) c1470153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470153));
	wire w1540153;
	torch #(1'b0) c1540153 (.i_clk(tick), .i_in(), .o_out(w1540153));
	wire w1580153;
	torch #(1'b0) c1580153 (.i_clk(tick), .i_in(), .o_out(w1580153));
	wire w1620153;
	torch #(1'b0) c1620153 (.i_clk(tick), .i_in(), .o_out(w1620153));
	wire w1660153;
	torch #(1'b0) c1660153 (.i_clk(tick), .i_in(), .o_out(w1660153));
	wire w1700153;
	torch #(1'b0) c1700153 (.i_clk(tick), .i_in(), .o_out(w1700153));
	wire w1740153;
	torch #(1'b0) c1740153 (.i_clk(tick), .i_in(), .o_out(w1740153));
	wire w1780153;
	torch #(1'b0) c1780153 (.i_clk(tick), .i_in(), .o_out(w1780153));
	wire w1470154;
	repeater #(1, 1'b0, 0, 0) c1470154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470154));
	wire w1470155;
	repeater #(1, 1'b0, 0, 0) c1470155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470155));
	wire w1540158;

	wire w1580158;

	wire w1620158;

	wire w1660158;

	wire w1700158;

	wire w1740158;

	wire w1780158;

	wire w1550167;
	torch #(1'b1) c1550167 (.i_clk(tick), .i_in(), .o_out(w1550167));
	wire w1590167;
	torch #(1'b1) c1590167 (.i_clk(tick), .i_in(), .o_out(w1590167));
	wire w1630167;
	torch #(1'b1) c1630167 (.i_clk(tick), .i_in(), .o_out(w1630167));
	wire w1670167;
	torch #(1'b1) c1670167 (.i_clk(tick), .i_in(), .o_out(w1670167));
	wire w1710167;
	torch #(1'b1) c1710167 (.i_clk(tick), .i_in(), .o_out(w1710167));
	wire w1750167;
	torch #(1'b1) c1750167 (.i_clk(tick), .i_in(), .o_out(w1750167));
	wire w1790167;
	torch #(1'b1) c1790167 (.i_clk(tick), .i_in(), .o_out(w1790167));
	wire w1540169;
	torch #(1'b0) c1540169 (.i_clk(tick), .i_in(), .o_out(w1540169));
	wire w1580169;
	torch #(1'b0) c1580169 (.i_clk(tick), .i_in(), .o_out(w1580169));
	wire w1620169;
	torch #(1'b0) c1620169 (.i_clk(tick), .i_in(), .o_out(w1620169));
	wire w1660169;
	torch #(1'b0) c1660169 (.i_clk(tick), .i_in(), .o_out(w1660169));
	wire w1700169;
	torch #(1'b0) c1700169 (.i_clk(tick), .i_in(), .o_out(w1700169));
	wire w1740169;
	torch #(1'b0) c1740169 (.i_clk(tick), .i_in(), .o_out(w1740169));
	wire w1780169;
	torch #(1'b0) c1780169 (.i_clk(tick), .i_in(), .o_out(w1780169));
	wire w1520172;
	assign outputs[96] = ();
	wire w1540172;
	assign outputs[97] = ();
	wire w1560172;
	assign outputs[98] = ();
	wire w1580172;
	assign outputs[99] = ();
	wire w1600172;
	assign outputs[100] = ();
	wire w1620172;
	assign outputs[101] = ();
	wire w1640172;
	assign outputs[102] = ();
	wire w1660172;
	assign outputs[103] = ();
	wire w1680172;
	assign outputs[104] = ();
	wire w1700172;
	assign outputs[105] = ();
	wire w1720172;
	assign outputs[106] = ();
	wire w1740172;
	assign outputs[107] = ();
	wire w1760172;
	assign outputs[108] = ();
	wire w1780172;
	assign outputs[109] = ();
	wire w1520173;
	repeater #(1, 1'b0, 0, 0) c1520173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520173));
	wire w1540173;
	repeater #(1, 1'b0, 0, 0) c1540173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1540173));
	wire w1560173;
	repeater #(1, 1'b0, 0, 0) c1560173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560173));
	wire w1580173;
	repeater #(1, 1'b0, 0, 0) c1580173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580173));
	wire w1600173;
	repeater #(1, 1'b0, 0, 0) c1600173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1600173));
	wire w1620173;
	repeater #(1, 1'b0, 0, 0) c1620173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1620173));
	wire w1640173;
	repeater #(1, 1'b0, 0, 0) c1640173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640173));
	wire w1660173;
	repeater #(1, 1'b0, 0, 0) c1660173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1660173));
	wire w1680173;
	repeater #(1, 1'b0, 0, 0) c1680173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1680173));
	wire w1700173;
	repeater #(1, 1'b0, 0, 0) c1700173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1700173));
	wire w1720173;
	repeater #(1, 1'b0, 0, 0) c1720173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1720173));
	wire w1740173;
	repeater #(1, 1'b0, 0, 0) c1740173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1740173));
	wire w1760173;
	repeater #(1, 1'b0, 0, 0) c1760173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1760173));
	wire w1780173;
	repeater #(1, 1'b0, 0, 0) c1780173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1780173));
	wire w15311;
	repeater #(2, 1'b1, 0, 0) c15311 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15311));
	wire w15711;
	repeater #(2, 1'b1, 0, 0) c15711 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15711));
	wire w16111;
	repeater #(2, 1'b1, 0, 0) c16111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16111));
	wire w16511;
	repeater #(2, 1'b1, 0, 0) c16511 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16511));
	wire w16911;
	repeater #(2, 1'b1, 0, 0) c16911 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16911));
	wire w17311;
	repeater #(2, 1'b1, 0, 0) c17311 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17311));
	wire w17711;
	repeater #(2, 1'b1, 0, 0) c17711 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17711));
	wire w15116;
	repeater #(1, 1'b1, 0, 0) c15116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15116));
	wire w15516;
	repeater #(1, 1'b1, 0, 0) c15516 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15516));
	wire w15916;
	repeater #(1, 1'b1, 0, 0) c15916 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15916));
	wire w16316;
	repeater #(1, 1'b1, 0, 0) c16316 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16316));
	wire w16716;
	repeater #(1, 1'b1, 0, 0) c16716 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16716));
	wire w17116;
	repeater #(1, 1'b1, 0, 0) c17116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17116));
	wire w17516;
	repeater #(1, 1'b1, 0, 0) c17516 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17516));
	wire w15317;

	wire w15717;

	wire w16117;

	wire w16517;

	wire w16917;

	wire w17317;

	wire w17717;

	wire w15218;

	wire w15618;

	wire w16018;

	wire w16418;

	wire w16818;

	wire w17218;

	wire w17618;

	wire w15319;
	torch #(1'b1) c15319 (.i_clk(tick), .i_in(), .o_out(w15319));
	wire w15719;
	torch #(1'b1) c15719 (.i_clk(tick), .i_in(), .o_out(w15719));
	wire w16119;
	torch #(1'b1) c16119 (.i_clk(tick), .i_in(), .o_out(w16119));
	wire w16519;
	torch #(1'b1) c16519 (.i_clk(tick), .i_in(), .o_out(w16519));
	wire w16919;
	torch #(1'b1) c16919 (.i_clk(tick), .i_in(), .o_out(w16919));
	wire w17319;
	torch #(1'b1) c17319 (.i_clk(tick), .i_in(), .o_out(w17319));
	wire w17719;
	torch #(1'b1) c17719 (.i_clk(tick), .i_in(), .o_out(w17719));
	wire w151110;
	repeater #(1, 1'b1, 0, 0) c151110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151110));
	wire w155110;
	repeater #(1, 1'b1, 0, 0) c155110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155110));
	wire w159110;
	repeater #(1, 1'b1, 0, 0) c159110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159110));
	wire w163110;
	repeater #(1, 1'b1, 0, 0) c163110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163110));
	wire w167110;
	repeater #(1, 1'b1, 0, 0) c167110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167110));
	wire w171110;
	repeater #(1, 1'b1, 0, 0) c171110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171110));
	wire w175110;
	repeater #(1, 1'b1, 0, 0) c175110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175110));
	wire w179123;
	assign outputs[110] = ();
	wire w179125;
	assign outputs[111] = ();
	wire w179127;
	assign outputs[112] = ();
	wire w179129;
	assign outputs[113] = ();
	wire w185135;
	assign outputs[114] = ();
	wire w105143;
	repeater #(1, 1'b0, 0, 0) c105143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105143));
	wire w104144;
	torch #(1'b0) c104144 (.i_clk(tick), .i_in(), .o_out(w104144));
	wire w153182;
	torch #(1'b1) c153182 (.i_clk(tick), .i_in(), .o_out(w153182));
	wire w157182;
	torch #(1'b1) c157182 (.i_clk(tick), .i_in(), .o_out(w157182));
	wire w161182;
	torch #(1'b1) c161182 (.i_clk(tick), .i_in(), .o_out(w161182));
	wire w165182;
	torch #(1'b1) c165182 (.i_clk(tick), .i_in(), .o_out(w165182));
	wire w169182;
	torch #(1'b1) c169182 (.i_clk(tick), .i_in(), .o_out(w169182));
	wire w173182;
	torch #(1'b1) c173182 (.i_clk(tick), .i_in(), .o_out(w173182));
	wire w177182;
	torch #(1'b1) c177182 (.i_clk(tick), .i_in(), .o_out(w177182));
	wire w154185;
	repeater #(2, 1'b0, 0, 0) c154185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154185));
	wire w158185;
	repeater #(2, 1'b0, 0, 0) c158185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158185));
	wire w162185;
	repeater #(2, 1'b0, 0, 0) c162185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162185));
	wire w166185;
	repeater #(2, 1'b0, 0, 0) c166185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166185));
	wire w170185;
	repeater #(1, 1'b0, 0, 0) c170185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170185));
	wire w174185;
	repeater #(1, 1'b0, 0, 0) c174185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174185));
	wire w178185;
	repeater #(1, 1'b0, 0, 0) c178185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178185));
	wire w167186;
	repeater #(1, 1'b0, 0, 0) c167186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167186));
	wire w179186;
	repeater #(1, 1'b0, 0, 0) c179186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179186));
	wire w113199;
	repeater #(1, 1'b0, 0, 0) c113199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113199));
	wire w1541103;

	wire w1581103;

	wire w1621103;

	wire w1661103;

	wire w1701103;

	wire w1741103;

	wire w1781103;

	wire w1541104;
	repeater #(1, 1'b1, 0, 0) c1541104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541104));
	wire w1581104;
	repeater #(1, 1'b1, 0, 0) c1581104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581104));
	wire w1621104;
	repeater #(1, 1'b1, 0, 0) c1621104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621104));
	wire w1661104;
	repeater #(1, 1'b1, 0, 0) c1661104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661104));
	wire w1701104;
	repeater #(1, 1'b1, 0, 0) c1701104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701104));
	wire w1741104;
	repeater #(1, 1'b1, 0, 0) c1741104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741104));
	wire w1781104;
	repeater #(1, 1'b1, 0, 0) c1781104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781104));
	wire w1541119;

	wire w1581119;

	wire w1621119;

	wire w1661119;

	wire w1701119;

	wire w1741119;

	wire w1781119;

	wire w1541120;
	repeater #(1, 1'b1, 0, 0) c1541120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541120));
	wire w1581120;
	repeater #(1, 1'b1, 0, 0) c1581120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581120));
	wire w1621120;
	repeater #(1, 1'b1, 0, 0) c1621120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621120));
	wire w1661120;
	repeater #(1, 1'b1, 0, 0) c1661120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661120));
	wire w1701120;
	repeater #(1, 1'b1, 0, 0) c1701120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701120));
	wire w1741120;
	repeater #(1, 1'b1, 0, 0) c1741120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741120));
	wire w1781120;
	repeater #(1, 1'b1, 0, 0) c1781120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781120));
	wire w1541135;

	wire w1581135;

	wire w1621135;

	wire w1661135;

	wire w1701135;

	wire w1741135;

	wire w1781135;

	wire w13800;
	repeater #(1, 1'b1, 0, 0) c13800 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13800));
	wire w14200;
	repeater #(1, 1'b1, 0, 0) c14200 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14200));
	wire w14600;
	repeater #(1, 1'b1, 0, 0) c14600 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14600));
	wire w15000;
	repeater #(1, 1'b1, 0, 0) c15000 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15000));
	wire w15400;
	repeater #(1, 1'b1, 0, 0) c15400 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15400));
	wire w15800;
	repeater #(1, 1'b1, 0, 0) c15800 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15800));
	wire w16200;
	repeater #(1, 1'b1, 0, 0) c16200 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16200));
	wire w138015;

	wire w142015;

	wire w146015;

	wire w150015;

	wire w154015;

	wire w158015;

	wire w162015;

	wire w138016;
	repeater #(1, 1'b1, 0, 0) c138016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138016));
	wire w142016;
	repeater #(1, 1'b1, 0, 0) c142016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142016));
	wire w146016;
	repeater #(1, 1'b1, 0, 0) c146016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146016));
	wire w150016;
	repeater #(1, 1'b1, 0, 0) c150016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150016));
	wire w154016;
	repeater #(1, 1'b1, 0, 0) c154016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154016));
	wire w158016;
	repeater #(1, 1'b1, 0, 0) c158016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158016));
	wire w162016;
	repeater #(1, 1'b1, 0, 0) c162016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162016));
	wire w138031;

	wire w142031;

	wire w146031;

	wire w150031;

	wire w154031;

	wire w158031;

	wire w162031;

	wire w138032;
	repeater #(1, 1'b1, 0, 0) c138032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138032));
	wire w142032;
	repeater #(1, 1'b1, 0, 0) c142032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142032));
	wire w146032;
	repeater #(1, 1'b1, 0, 0) c146032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146032));
	wire w150032;
	repeater #(1, 1'b1, 0, 0) c150032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150032));
	wire w154032;
	repeater #(1, 1'b1, 0, 0) c154032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154032));
	wire w158032;
	repeater #(1, 1'b1, 0, 0) c158032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158032));
	wire w162032;
	repeater #(1, 1'b1, 0, 0) c162032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162032));
	wire w137040;
	torch #(1'b1) c137040 (.i_clk(tick), .i_in(), .o_out(w137040));
	wire w141040;
	torch #(1'b1) c141040 (.i_clk(tick), .i_in(), .o_out(w141040));
	wire w145040;
	torch #(1'b1) c145040 (.i_clk(tick), .i_in(), .o_out(w145040));
	wire w149040;
	torch #(1'b1) c149040 (.i_clk(tick), .i_in(), .o_out(w149040));
	wire w153040;
	torch #(1'b1) c153040 (.i_clk(tick), .i_in(), .o_out(w153040));
	wire w157040;
	torch #(1'b1) c157040 (.i_clk(tick), .i_in(), .o_out(w157040));
	wire w161040;
	torch #(1'b1) c161040 (.i_clk(tick), .i_in(), .o_out(w161040));
	wire w137044;
	torch #(1'b1) c137044 (.i_clk(tick), .i_in(), .o_out(w137044));
	wire w141044;
	torch #(1'b1) c141044 (.i_clk(tick), .i_in(), .o_out(w141044));
	wire w145044;
	torch #(1'b1) c145044 (.i_clk(tick), .i_in(), .o_out(w145044));
	wire w149044;
	torch #(1'b1) c149044 (.i_clk(tick), .i_in(), .o_out(w149044));
	wire w153044;
	torch #(1'b1) c153044 (.i_clk(tick), .i_in(), .o_out(w153044));
	wire w157044;
	torch #(1'b1) c157044 (.i_clk(tick), .i_in(), .o_out(w157044));
	wire w161044;
	torch #(1'b1) c161044 (.i_clk(tick), .i_in(), .o_out(w161044));
	wire w136052;
	torch #(1'b1) c136052 (.i_clk(tick), .i_in(), .o_out(w136052));
	wire w140052;
	torch #(1'b1) c140052 (.i_clk(tick), .i_in(), .o_out(w140052));
	wire w144052;
	torch #(1'b1) c144052 (.i_clk(tick), .i_in(), .o_out(w144052));
	wire w148052;
	torch #(1'b1) c148052 (.i_clk(tick), .i_in(), .o_out(w148052));
	wire w152052;
	torch #(1'b1) c152052 (.i_clk(tick), .i_in(), .o_out(w152052));
	wire w156052;
	torch #(1'b1) c156052 (.i_clk(tick), .i_in(), .o_out(w156052));
	wire w160052;
	torch #(1'b1) c160052 (.i_clk(tick), .i_in(), .o_out(w160052));
	wire w148066;
	repeater #(1, 1'b0, 0, 0) c148066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148066));
	wire w163066;
	repeater #(1, 1'b0, 0, 0) c163066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163066));
	wire w148068;
	repeater #(1, 1'b0, 0, 0) c148068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148068));
	wire w163068;
	repeater #(1, 1'b0, 0, 0) c163068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163068));
	wire w167068;
	repeater #(1, 1'b0, 0, 0) c167068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167068));
	wire w148070;
	repeater #(1, 1'b0, 0, 0) c148070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148070));
	wire w163070;
	repeater #(1, 1'b0, 0, 0) c163070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163070));
	wire w148072;
	repeater #(1, 1'b0, 0, 0) c148072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148072));
	wire w163072;
	repeater #(1, 1'b0, 0, 0) c163072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163072));
	wire w169074;
	repeater #(1, 1'b0, 0, 0) c169074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169074));
	wire w171074;

	wire w172074;
	repeater #(4, 1'b1, 0, 0) c172074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172074));
	wire w171075;
	repeater #(1, 1'b1, 0, 0) c171075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171075));
	wire w172076;
	repeater #(4, 1'b1, 0, 0) c172076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w172076));
	wire w89085;
	repeater #(1, 1'b0, 0, 0) c89085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89085));
	wire w88086;
	torch #(1'b0) c88086 (.i_clk(tick), .i_in(), .o_out(w88086));
	wire w1320129;
	torch #(1'b0) c1320129 (.i_clk(tick), .i_in(), .o_out(w1320129));
	wire w1310134;
	repeater #(1, 1'b0, 0, 0) c1310134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310134));
	wire w1420135;
	repeater #(1, 1'b0, 0, 0) c1420135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420135));
	wire w1610135;
	repeater #(1, 1'b0, 0, 0) c1610135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610135));
	wire w1490136;
	repeater #(1, 1'b0, 0, 0) c1490136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490136));
	wire w1340137;
	repeater #(1, 1'b0, 0, 0) c1340137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340137));
	wire w1360137;

	wire w980141;

	wire w1340143;
	repeater #(1, 1'b0, 0, 0) c1340143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340143));
	wire w1360143;

	wire w1370143;
	repeater #(1, 1'b0, 0, 0) c1370143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370143));
	wire w1460143;
	repeater #(1, 1'b0, 0, 0) c1460143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460143));
	wire w1470143;
	repeater #(1, 1'b0, 0, 0) c1470143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470143));
	wire w1480143;
	repeater #(1, 1'b0, 0, 0) c1480143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1480143));
	wire w1490144;
	repeater #(1, 1'b0, 0, 0) c1490144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490144));
	wire w1310148;
	repeater #(1, 1'b0, 0, 0) c1310148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310148));
	wire w1310149;
	repeater #(1, 1'b0, 0, 0) c1310149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310149));
	wire w1310150;
	repeater #(1, 1'b0, 0, 0) c1310150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310150));
	wire w1420151;
	repeater #(1, 1'b0, 0, 0) c1420151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420151));
	wire w1610151;
	repeater #(1, 1'b0, 0, 0) c1610151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610151));
	wire w1490152;
	repeater #(1, 1'b0, 0, 0) c1490152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490152));
	wire w1340153;
	repeater #(1, 1'b0, 0, 0) c1340153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340153));
	wire w1360153;

	wire w1340159;
	repeater #(1, 1'b0, 0, 0) c1340159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340159));
	wire w1360159;

	wire w1370159;
	repeater #(1, 1'b0, 0, 0) c1370159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370159));
	wire w1460159;
	repeater #(1, 1'b0, 0, 0) c1460159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460159));
	wire w1470159;
	repeater #(1, 1'b0, 0, 0) c1470159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470159));
	wire w1480159;
	repeater #(1, 1'b0, 0, 0) c1480159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1480159));
	wire w1490160;
	repeater #(1, 1'b0, 0, 0) c1490160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490160));
	wire w1310164;
	repeater #(1, 1'b0, 0, 0) c1310164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310164));
	wire w1310165;
	repeater #(1, 1'b0, 0, 0) c1310165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310165));
	wire w1310166;
	repeater #(1, 1'b0, 0, 0) c1310166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1310166));
	wire w1420167;
	repeater #(1, 1'b0, 0, 0) c1420167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420167));
	wire w1610167;
	repeater #(1, 1'b0, 0, 0) c1610167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610167));
	wire w1490168;
	repeater #(1, 1'b0, 0, 0) c1490168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490168));
	wire w1340169;
	repeater #(1, 1'b0, 0, 0) c1340169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340169));
	wire w1360169;

	wire w1340175;
	repeater #(1, 1'b0, 0, 0) c1340175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340175));
	wire w1360175;

	wire w1370175;
	repeater #(1, 1'b0, 0, 0) c1370175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370175));
	wire w1460175;
	repeater #(1, 1'b0, 0, 0) c1460175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460175));
	wire w1470175;
	repeater #(1, 1'b0, 0, 0) c1470175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470175));
	wire w1480175;
	repeater #(1, 1'b0, 0, 0) c1480175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1480175));
	wire w1360176;
	repeater #(1, 1'b0, 0, 0) c1360176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1360176));
	wire w1490176;
	repeater #(1, 1'b0, 0, 0) c1490176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1490176));
	wire w13111;
	repeater #(1, 1'b0, 0, 0) c13111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13111));
	wire w13112;
	repeater #(1, 1'b0, 0, 0) c13112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13112));
	wire w13113;
	repeater #(1, 1'b0, 0, 0) c13113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13113));
	wire w14214;
	repeater #(1, 1'b0, 0, 0) c14214 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14214));
	wire w16114;
	repeater #(1, 1'b0, 0, 0) c16114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16114));
	wire w14915;
	repeater #(1, 1'b0, 0, 0) c14915 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14915));
	wire w13416;
	repeater #(1, 1'b0, 0, 0) c13416 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13416));
	wire w13616;

	wire w134112;
	repeater #(1, 1'b0, 0, 0) c134112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134112));
	wire w136112;

	wire w137112;
	repeater #(1, 1'b0, 0, 0) c137112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137112));
	wire w146112;
	repeater #(1, 1'b0, 0, 0) c146112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146112));
	wire w147112;
	repeater #(1, 1'b0, 0, 0) c147112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147112));
	wire w148112;
	repeater #(1, 1'b0, 0, 0) c148112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148112));
	wire w149113;
	repeater #(1, 1'b0, 0, 0) c149113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149113));
	wire w131117;
	repeater #(1, 1'b0, 0, 0) c131117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131117));
	wire w131118;
	repeater #(1, 1'b0, 0, 0) c131118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131118));
	wire w131119;
	repeater #(1, 1'b0, 0, 0) c131119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131119));
	wire w142120;
	repeater #(1, 1'b0, 0, 0) c142120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142120));
	wire w161120;
	repeater #(1, 1'b0, 0, 0) c161120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161120));
	wire w149121;
	repeater #(1, 1'b0, 0, 0) c149121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149121));
	wire w134122;
	repeater #(1, 1'b0, 0, 0) c134122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134122));
	wire w136122;

	wire w134128;
	repeater #(1, 1'b0, 0, 0) c134128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134128));
	wire w136128;

	wire w137128;
	repeater #(1, 1'b0, 0, 0) c137128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w137128));
	wire w146128;
	repeater #(1, 1'b0, 0, 0) c146128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146128));
	wire w147128;
	repeater #(1, 1'b0, 0, 0) c147128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147128));
	wire w148128;
	repeater #(1, 1'b0, 0, 0) c148128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148128));
	wire w149129;
	repeater #(1, 1'b0, 0, 0) c149129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149129));
	wire w135143;
	repeater #(1, 1'b0, 0, 0) c135143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135143));
	wire w139143;
	repeater #(1, 1'b0, 0, 0) c139143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139143));
	wire w143143;
	repeater #(1, 1'b0, 0, 0) c143143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143143));
	wire w147143;
	repeater #(1, 1'b0, 0, 0) c147143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147143));
	wire w151143;
	repeater #(1, 1'b0, 0, 0) c151143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151143));
	wire w155143;
	repeater #(1, 1'b0, 0, 0) c155143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155143));
	wire w159143;
	repeater #(1, 1'b0, 0, 0) c159143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159143));
	wire w136145;

	wire w140145;

	wire w144145;

	wire w148145;

	wire w152145;

	wire w156145;

	wire w160145;

	wire w136146;

	wire w140146;

	wire w144146;

	wire w148146;

	wire w152146;

	wire w156146;

	wire w160146;

	wire w135149;
	repeater #(1, 1'b1, 0, 0) c135149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135149));
	wire w139149;
	repeater #(1, 1'b1, 0, 0) c139149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139149));
	wire w143149;
	repeater #(1, 1'b1, 0, 0) c143149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143149));
	wire w147149;
	repeater #(1, 1'b1, 0, 0) c147149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147149));
	wire w151149;
	repeater #(1, 1'b1, 0, 0) c151149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151149));
	wire w155149;
	repeater #(1, 1'b1, 0, 0) c155149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155149));
	wire w159149;
	repeater #(1, 1'b1, 0, 0) c159149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159149));
	wire w137150;

	wire w141150;

	wire w145150;

	wire w149150;

	wire w153150;

	wire w157150;

	wire w161150;

	wire w136151;

	wire w140151;

	wire w144151;

	wire w148151;

	wire w152151;

	wire w156151;

	wire w160151;

	wire w139166;
	torch #(1'b1) c139166 (.i_clk(tick), .i_in(), .o_out(w139166));
	wire w145166;
	torch #(1'b1) c145166 (.i_clk(tick), .i_in(), .o_out(w145166));
	wire w153166;
	torch #(1'b1) c153166 (.i_clk(tick), .i_in(), .o_out(w153166));
	wire w161166;
	torch #(1'b1) c161166 (.i_clk(tick), .i_in(), .o_out(w161166));
	wire w139168;
	torch #(1'b1) c139168 (.i_clk(tick), .i_in(), .o_out(w139168));
	wire w141168;
	torch #(1'b1) c141168 (.i_clk(tick), .i_in(), .o_out(w141168));
	wire w153168;
	torch #(1'b1) c153168 (.i_clk(tick), .i_in(), .o_out(w153168));
	wire w157168;
	torch #(1'b1) c157168 (.i_clk(tick), .i_in(), .o_out(w157168));
	wire w139170;
	torch #(1'b1) c139170 (.i_clk(tick), .i_in(), .o_out(w139170));
	wire w141170;
	torch #(1'b1) c141170 (.i_clk(tick), .i_in(), .o_out(w141170));
	wire w145170;
	torch #(1'b1) c145170 (.i_clk(tick), .i_in(), .o_out(w145170));
	wire w149170;
	torch #(1'b1) c149170 (.i_clk(tick), .i_in(), .o_out(w149170));
	wire w139172;
	torch #(1'b1) c139172 (.i_clk(tick), .i_in(), .o_out(w139172));
	wire w141172;
	torch #(1'b1) c141172 (.i_clk(tick), .i_in(), .o_out(w141172));
	wire w145172;
	torch #(1'b1) c145172 (.i_clk(tick), .i_in(), .o_out(w145172));
	wire w149172;
	torch #(1'b1) c149172 (.i_clk(tick), .i_in(), .o_out(w149172));
	wire w153172;
	torch #(1'b1) c153172 (.i_clk(tick), .i_in(), .o_out(w153172));
	wire w157172;
	torch #(1'b1) c157172 (.i_clk(tick), .i_in(), .o_out(w157172));
	wire w161172;
	torch #(1'b1) c161172 (.i_clk(tick), .i_in(), .o_out(w161172));
	wire w169178;
	assign outputs[115] = ();
	wire w89187;
	repeater #(1, 1'b0, 0, 0) c89187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89187));
	wire w1291116;
	repeater #(1, 1'b0, 0, 0) c1291116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1291116));
	wire w1291126;
	repeater #(1, 1'b0, 0, 0) c1291126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1291126));
	wire w1311128;

	wire w1331128;

	wire w8206;
	repeater #(1, 1'b1, 0, 0) c8206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8206));
	wire w122093;
	torch #(1'b1) c122093 (.i_clk(tick), .i_in(), .o_out(w122093));
	wire w126093;
	torch #(1'b1) c126093 (.i_clk(tick), .i_in(), .o_out(w126093));
	wire w130093;
	torch #(1'b1) c130093 (.i_clk(tick), .i_in(), .o_out(w130093));
	wire w134093;
	torch #(1'b1) c134093 (.i_clk(tick), .i_in(), .o_out(w134093));
	wire w138093;
	torch #(1'b1) c138093 (.i_clk(tick), .i_in(), .o_out(w138093));
	wire w142093;
	torch #(1'b1) c142093 (.i_clk(tick), .i_in(), .o_out(w142093));
	wire w146093;
	torch #(1'b1) c146093 (.i_clk(tick), .i_in(), .o_out(w146093));
	wire w1220108;
	torch #(1'b0) c1220108 (.i_clk(tick), .i_in(), .o_out(w1220108));
	wire w1260108;
	torch #(1'b0) c1260108 (.i_clk(tick), .i_in(), .o_out(w1260108));
	wire w1300108;
	torch #(1'b0) c1300108 (.i_clk(tick), .i_in(), .o_out(w1300108));
	wire w1340108;
	torch #(1'b0) c1340108 (.i_clk(tick), .i_in(), .o_out(w1340108));
	wire w1380108;
	torch #(1'b0) c1380108 (.i_clk(tick), .i_in(), .o_out(w1380108));
	wire w1420108;
	torch #(1'b0) c1420108 (.i_clk(tick), .i_in(), .o_out(w1420108));
	wire w1460108;
	torch #(1'b0) c1460108 (.i_clk(tick), .i_in(), .o_out(w1460108));
	wire w1530117;
	repeater #(1, 1'b0, 0, 0) c1530117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1530117));
	wire w1550117;

	wire w1560117;
	repeater #(4, 1'b0, 0, 0) c1560117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560117));
	wire w1550118;
	repeater #(1, 1'b0, 0, 0) c1550118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550118));
	wire w1560119;
	repeater #(4, 1'b0, 0, 0) c1560119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1560119));
	wire w1100158;
	repeater #(1, 1'b0, 0, 0) c1100158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1100158));
	wire w1190168;
	repeater #(1, 1'b0, 0, 0) c1190168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190168));
	wire w1190169;
	repeater #(2, 1'b0, 0, 0) c1190169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190169));
	wire w1190170;
	repeater #(2, 1'b0, 0, 0) c1190170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190170));
	wire w1190171;
	repeater #(2, 1'b0, 0, 0) c1190171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190171));
	wire w1190172;
	repeater #(2, 1'b0, 0, 0) c1190172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1190172));
	wire w1150178;
	repeater #(1, 1'b0, 0, 0) c1150178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1150178));
	wire w8115;

	wire w120111;
	repeater #(1, 1'b0, 0, 0) c120111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120111));
	wire w115112;
	repeater #(1, 1'b0, 0, 0) c115112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115112));
	wire w120112;
	repeater #(1, 1'b0, 0, 0) c120112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120112));
	wire w115113;
	repeater #(1, 1'b0, 0, 0) c115113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115113));
	wire w115114;
	repeater #(1, 1'b0, 0, 0) c115114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115114));
	wire w120116;
	repeater #(1, 1'b0, 0, 0) c120116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120116));
	wire w120127;
	repeater #(1, 1'b0, 0, 0) c120127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120127));
	wire w115128;
	repeater #(1, 1'b0, 0, 0) c115128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115128));
	wire w120128;
	repeater #(1, 1'b0, 0, 0) c120128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120128));
	wire w115129;
	repeater #(1, 1'b0, 0, 0) c115129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115129));
	wire w115130;
	repeater #(1, 1'b0, 0, 0) c115130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115130));
	wire w124130;
	repeater #(1, 1'b0, 0, 0) c124130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124130));
	wire w128130;
	repeater #(1, 1'b0, 0, 0) c128130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128130));
	wire w132130;
	repeater #(1, 1'b0, 0, 0) c132130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132130));
	wire w136130;
	repeater #(1, 1'b0, 0, 0) c136130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136130));
	wire w140130;
	repeater #(1, 1'b0, 0, 0) c140130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140130));
	wire w144130;
	repeater #(1, 1'b0, 0, 0) c144130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144130));
	wire w148130;
	repeater #(1, 1'b0, 0, 0) c148130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148130));
	wire w124131;
	repeater #(4, 1'b0, 0, 0) c124131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124131));
	wire w128131;
	repeater #(4, 1'b0, 0, 0) c128131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128131));
	wire w132131;
	repeater #(4, 1'b0, 0, 0) c132131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132131));
	wire w136131;
	repeater #(4, 1'b0, 0, 0) c136131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136131));
	wire w140131;
	repeater #(4, 1'b0, 0, 0) c140131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140131));
	wire w144131;
	repeater #(4, 1'b0, 0, 0) c144131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144131));
	wire w148131;
	repeater #(4, 1'b0, 0, 0) c148131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148131));
	wire w120132;
	repeater #(1, 1'b0, 0, 0) c120132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120132));
	wire w120143;
	repeater #(1, 1'b0, 0, 0) c120143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120143));
	wire w115144;
	repeater #(1, 1'b0, 0, 0) c115144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115144));
	wire w120144;
	repeater #(1, 1'b0, 0, 0) c120144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120144));
	wire w115145;
	repeater #(1, 1'b0, 0, 0) c115145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115145));
	wire w115146;
	repeater #(1, 1'b0, 0, 0) c115146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115146));
	wire w124146;
	repeater #(3, 1'b0, 0, 0) c124146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124146));
	wire w128146;
	repeater #(3, 1'b0, 0, 0) c128146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128146));
	wire w132146;
	repeater #(3, 1'b0, 0, 0) c132146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132146));
	wire w136146;
	repeater #(3, 1'b0, 0, 0) c136146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136146));
	wire w140146;
	repeater #(3, 1'b0, 0, 0) c140146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140146));
	wire w144146;
	repeater #(3, 1'b0, 0, 0) c144146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144146));
	wire w148146;
	repeater #(3, 1'b0, 0, 0) c148146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148146));
	wire w124147;
	repeater #(4, 1'b0, 0, 0) c124147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124147));
	wire w128147;
	repeater #(4, 1'b0, 0, 0) c128147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128147));
	wire w132147;
	repeater #(4, 1'b0, 0, 0) c132147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132147));
	wire w136147;
	repeater #(4, 1'b0, 0, 0) c136147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136147));
	wire w140147;
	repeater #(4, 1'b0, 0, 0) c140147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140147));
	wire w144147;
	repeater #(4, 1'b0, 0, 0) c144147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144147));
	wire w148147;
	repeater #(4, 1'b0, 0, 0) c148147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148147));
	wire w120148;
	repeater #(1, 1'b0, 0, 0) c120148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120148));
	wire w124148;
	repeater #(4, 1'b0, 0, 0) c124148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124148));
	wire w128148;
	repeater #(4, 1'b0, 0, 0) c128148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128148));
	wire w132148;
	repeater #(4, 1'b0, 0, 0) c132148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132148));
	wire w136148;
	repeater #(4, 1'b0, 0, 0) c136148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136148));
	wire w140148;
	repeater #(4, 1'b0, 0, 0) c140148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140148));
	wire w144148;
	repeater #(4, 1'b0, 0, 0) c144148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144148));
	wire w148148;
	repeater #(4, 1'b0, 0, 0) c148148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148148));
	wire w124149;
	repeater #(4, 1'b0, 0, 0) c124149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124149));
	wire w128149;
	repeater #(4, 1'b0, 0, 0) c128149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128149));
	wire w132149;
	repeater #(4, 1'b0, 0, 0) c132149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132149));
	wire w136149;
	repeater #(4, 1'b0, 0, 0) c136149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136149));
	wire w140149;
	repeater #(4, 1'b0, 0, 0) c140149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140149));
	wire w144149;
	repeater #(4, 1'b0, 0, 0) c144149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144149));
	wire w148149;
	repeater #(4, 1'b0, 0, 0) c148149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148149));
	wire w124150;
	repeater #(4, 1'b0, 0, 0) c124150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124150));
	wire w128150;
	repeater #(4, 1'b0, 0, 0) c128150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128150));
	wire w132150;
	repeater #(4, 1'b0, 0, 0) c132150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132150));
	wire w136150;
	repeater #(4, 1'b0, 0, 0) c136150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136150));
	wire w140150;
	repeater #(4, 1'b0, 0, 0) c140150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140150));
	wire w144150;
	repeater #(4, 1'b0, 0, 0) c144150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144150));
	wire w148150;
	repeater #(4, 1'b0, 0, 0) c148150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148150));
	wire w124151;
	repeater #(4, 1'b0, 0, 0) c124151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124151));
	wire w128151;
	repeater #(4, 1'b0, 0, 0) c128151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128151));
	wire w132151;
	repeater #(4, 1'b0, 0, 0) c132151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132151));
	wire w136151;
	repeater #(4, 1'b0, 0, 0) c136151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136151));
	wire w140151;
	repeater #(4, 1'b0, 0, 0) c140151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140151));
	wire w144151;
	repeater #(4, 1'b0, 0, 0) c144151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144151));
	wire w148151;
	repeater #(4, 1'b0, 0, 0) c148151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148151));
	wire w124152;
	repeater #(4, 1'b0, 0, 0) c124152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124152));
	wire w128152;
	repeater #(4, 1'b0, 0, 0) c128152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128152));
	wire w132152;
	repeater #(4, 1'b0, 0, 0) c132152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132152));
	wire w136152;
	repeater #(4, 1'b0, 0, 0) c136152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136152));
	wire w140152;
	repeater #(4, 1'b0, 0, 0) c140152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140152));
	wire w144152;
	repeater #(4, 1'b0, 0, 0) c144152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144152));
	wire w148152;
	repeater #(4, 1'b0, 0, 0) c148152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148152));
	wire w124153;
	repeater #(4, 1'b0, 0, 0) c124153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124153));
	wire w128153;
	repeater #(4, 1'b0, 0, 0) c128153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128153));
	wire w132153;
	repeater #(4, 1'b0, 0, 0) c132153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132153));
	wire w136153;
	repeater #(4, 1'b0, 0, 0) c136153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136153));
	wire w140153;
	repeater #(4, 1'b0, 0, 0) c140153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140153));
	wire w144153;
	repeater #(4, 1'b0, 0, 0) c144153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144153));
	wire w148153;
	repeater #(4, 1'b0, 0, 0) c148153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148153));
	wire w124154;
	repeater #(4, 1'b0, 0, 0) c124154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124154));
	wire w128154;
	repeater #(4, 1'b0, 0, 0) c128154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128154));
	wire w132154;
	repeater #(4, 1'b0, 0, 0) c132154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132154));
	wire w136154;
	repeater #(4, 1'b0, 0, 0) c136154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136154));
	wire w140154;
	repeater #(4, 1'b0, 0, 0) c140154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140154));
	wire w144154;
	repeater #(4, 1'b0, 0, 0) c144154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144154));
	wire w148154;
	repeater #(4, 1'b0, 0, 0) c148154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148154));
	wire w120159;
	repeater #(1, 1'b0, 0, 0) c120159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120159));
	wire w115160;
	repeater #(1, 1'b0, 0, 0) c115160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115160));
	wire w120160;
	repeater #(1, 1'b0, 0, 0) c120160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120160));
	wire w124160;
	repeater #(3, 1'b0, 0, 0) c124160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124160));
	wire w128160;
	repeater #(3, 1'b0, 0, 0) c128160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128160));
	wire w132160;
	repeater #(3, 1'b0, 0, 0) c132160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132160));
	wire w136160;
	repeater #(3, 1'b0, 0, 0) c136160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136160));
	wire w140160;
	repeater #(3, 1'b0, 0, 0) c140160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140160));
	wire w144160;
	repeater #(3, 1'b0, 0, 0) c144160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144160));
	wire w148160;
	repeater #(3, 1'b0, 0, 0) c148160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148160));
	wire w115161;
	repeater #(1, 1'b0, 0, 0) c115161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115161));
	wire w124161;
	repeater #(4, 1'b0, 0, 0) c124161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124161));
	wire w128161;
	repeater #(4, 1'b0, 0, 0) c128161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128161));
	wire w132161;
	repeater #(4, 1'b0, 0, 0) c132161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132161));
	wire w136161;
	repeater #(4, 1'b0, 0, 0) c136161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136161));
	wire w140161;
	repeater #(4, 1'b0, 0, 0) c140161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140161));
	wire w144161;
	repeater #(4, 1'b0, 0, 0) c144161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144161));
	wire w148161;
	repeater #(4, 1'b0, 0, 0) c148161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148161));
	wire w115162;
	repeater #(1, 1'b0, 0, 0) c115162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115162));
	wire w124162;
	repeater #(4, 1'b0, 0, 0) c124162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124162));
	wire w128162;
	repeater #(4, 1'b0, 0, 0) c128162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128162));
	wire w132162;
	repeater #(4, 1'b0, 0, 0) c132162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132162));
	wire w136162;
	repeater #(4, 1'b0, 0, 0) c136162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136162));
	wire w140162;
	repeater #(4, 1'b0, 0, 0) c140162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140162));
	wire w144162;
	repeater #(4, 1'b0, 0, 0) c144162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144162));
	wire w148162;
	repeater #(4, 1'b0, 0, 0) c148162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148162));
	wire w124163;
	repeater #(4, 1'b0, 0, 0) c124163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124163));
	wire w128163;
	repeater #(4, 1'b0, 0, 0) c128163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128163));
	wire w132163;
	repeater #(4, 1'b0, 0, 0) c132163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132163));
	wire w136163;
	repeater #(4, 1'b0, 0, 0) c136163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136163));
	wire w140163;
	repeater #(4, 1'b0, 0, 0) c140163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140163));
	wire w144163;
	repeater #(4, 1'b0, 0, 0) c144163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144163));
	wire w148163;
	repeater #(4, 1'b0, 0, 0) c148163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148163));
	wire w120164;
	repeater #(1, 1'b0, 0, 0) c120164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120164));
	wire w124164;
	repeater #(4, 1'b0, 0, 0) c124164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124164));
	wire w128164;
	repeater #(4, 1'b0, 0, 0) c128164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128164));
	wire w132164;
	repeater #(4, 1'b0, 0, 0) c132164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132164));
	wire w136164;
	repeater #(4, 1'b0, 0, 0) c136164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136164));
	wire w140164;
	repeater #(4, 1'b0, 0, 0) c140164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140164));
	wire w144164;
	repeater #(4, 1'b0, 0, 0) c144164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144164));
	wire w148164;
	repeater #(4, 1'b0, 0, 0) c148164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148164));
	wire w124165;
	repeater #(4, 1'b0, 0, 0) c124165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124165));
	wire w128165;
	repeater #(4, 1'b0, 0, 0) c128165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128165));
	wire w132165;
	repeater #(4, 1'b0, 0, 0) c132165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132165));
	wire w136165;
	repeater #(4, 1'b0, 0, 0) c136165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136165));
	wire w140165;
	repeater #(4, 1'b0, 0, 0) c140165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140165));
	wire w144165;
	repeater #(4, 1'b0, 0, 0) c144165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144165));
	wire w148165;
	repeater #(4, 1'b0, 0, 0) c148165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148165));
	wire w124166;
	repeater #(4, 1'b0, 0, 0) c124166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124166));
	wire w128166;
	repeater #(4, 1'b0, 0, 0) c128166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128166));
	wire w132166;
	repeater #(4, 1'b0, 0, 0) c132166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132166));
	wire w136166;
	repeater #(4, 1'b0, 0, 0) c136166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136166));
	wire w140166;
	repeater #(4, 1'b0, 0, 0) c140166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140166));
	wire w144166;
	repeater #(4, 1'b0, 0, 0) c144166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144166));
	wire w148166;
	repeater #(4, 1'b0, 0, 0) c148166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148166));
	wire w124167;
	repeater #(4, 1'b0, 0, 0) c124167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124167));
	wire w128167;
	repeater #(4, 1'b0, 0, 0) c128167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128167));
	wire w132167;
	repeater #(4, 1'b0, 0, 0) c132167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132167));
	wire w136167;
	repeater #(4, 1'b0, 0, 0) c136167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136167));
	wire w140167;
	repeater #(4, 1'b0, 0, 0) c140167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140167));
	wire w144167;
	repeater #(4, 1'b0, 0, 0) c144167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144167));
	wire w148167;
	repeater #(4, 1'b0, 0, 0) c148167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148167));
	wire w124168;
	repeater #(4, 1'b0, 0, 0) c124168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124168));
	wire w128168;
	repeater #(4, 1'b0, 0, 0) c128168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128168));
	wire w132168;
	repeater #(4, 1'b0, 0, 0) c132168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132168));
	wire w136168;
	repeater #(4, 1'b0, 0, 0) c136168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136168));
	wire w140168;
	repeater #(4, 1'b0, 0, 0) c140168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140168));
	wire w144168;
	repeater #(4, 1'b0, 0, 0) c144168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144168));
	wire w148168;
	repeater #(4, 1'b0, 0, 0) c148168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148168));
	wire w124169;
	repeater #(4, 1'b0, 0, 0) c124169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124169));
	wire w128169;
	repeater #(4, 1'b0, 0, 0) c128169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128169));
	wire w132169;
	repeater #(4, 1'b0, 0, 0) c132169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132169));
	wire w136169;
	repeater #(4, 1'b0, 0, 0) c136169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136169));
	wire w140169;
	repeater #(4, 1'b0, 0, 0) c140169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140169));
	wire w144169;
	repeater #(4, 1'b0, 0, 0) c144169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144169));
	wire w148169;
	repeater #(4, 1'b0, 0, 0) c148169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148169));
	wire w124170;
	repeater #(4, 1'b0, 0, 0) c124170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124170));
	wire w128170;
	repeater #(4, 1'b0, 0, 0) c128170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128170));
	wire w132170;
	repeater #(4, 1'b0, 0, 0) c132170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132170));
	wire w136170;
	repeater #(4, 1'b0, 0, 0) c136170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136170));
	wire w140170;
	repeater #(4, 1'b0, 0, 0) c140170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140170));
	wire w144170;
	repeater #(4, 1'b0, 0, 0) c144170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144170));
	wire w148170;
	repeater #(4, 1'b0, 0, 0) c148170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148170));
	wire w124171;
	repeater #(4, 1'b0, 0, 0) c124171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124171));
	wire w128171;
	repeater #(4, 1'b0, 0, 0) c128171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128171));
	wire w132171;
	repeater #(4, 1'b0, 0, 0) c132171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132171));
	wire w136171;
	repeater #(4, 1'b0, 0, 0) c136171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136171));
	wire w140171;
	repeater #(4, 1'b0, 0, 0) c140171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140171));
	wire w144171;
	repeater #(4, 1'b0, 0, 0) c144171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144171));
	wire w148171;
	repeater #(4, 1'b0, 0, 0) c148171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148171));
	wire w124172;
	repeater #(4, 1'b0, 0, 0) c124172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124172));
	wire w128172;
	repeater #(4, 1'b0, 0, 0) c128172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128172));
	wire w132172;
	repeater #(4, 1'b0, 0, 0) c132172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132172));
	wire w136172;
	repeater #(4, 1'b0, 0, 0) c136172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136172));
	wire w140172;
	repeater #(4, 1'b0, 0, 0) c140172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140172));
	wire w144172;
	repeater #(4, 1'b0, 0, 0) c144172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144172));
	wire w148172;
	repeater #(4, 1'b0, 0, 0) c148172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148172));
	wire w124173;
	repeater #(4, 1'b0, 0, 0) c124173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124173));
	wire w128173;
	repeater #(4, 1'b0, 0, 0) c128173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128173));
	wire w132173;
	repeater #(4, 1'b0, 0, 0) c132173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132173));
	wire w136173;
	repeater #(4, 1'b0, 0, 0) c136173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136173));
	wire w140173;
	repeater #(4, 1'b0, 0, 0) c140173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140173));
	wire w144173;
	repeater #(4, 1'b0, 0, 0) c144173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144173));
	wire w148173;
	repeater #(4, 1'b0, 0, 0) c148173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148173));
	wire w124174;
	repeater #(4, 1'b0, 0, 0) c124174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124174));
	wire w128174;
	repeater #(4, 1'b0, 0, 0) c128174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128174));
	wire w132174;
	repeater #(4, 1'b0, 0, 0) c132174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132174));
	wire w136174;
	repeater #(4, 1'b0, 0, 0) c136174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136174));
	wire w140174;
	repeater #(4, 1'b0, 0, 0) c140174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140174));
	wire w144174;
	repeater #(4, 1'b0, 0, 0) c144174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144174));
	wire w148174;
	repeater #(4, 1'b0, 0, 0) c148174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148174));
	wire w124175;
	repeater #(4, 1'b0, 0, 0) c124175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124175));
	wire w128175;
	repeater #(4, 1'b0, 0, 0) c128175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128175));
	wire w132175;
	repeater #(4, 1'b0, 0, 0) c132175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132175));
	wire w136175;
	repeater #(4, 1'b0, 0, 0) c136175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136175));
	wire w140175;
	repeater #(4, 1'b0, 0, 0) c140175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140175));
	wire w144175;
	repeater #(4, 1'b0, 0, 0) c144175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144175));
	wire w148175;
	repeater #(4, 1'b0, 0, 0) c148175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148175));
	wire w124176;
	repeater #(4, 1'b0, 0, 0) c124176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124176));
	wire w128176;
	repeater #(4, 1'b0, 0, 0) c128176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128176));
	wire w132176;
	repeater #(4, 1'b0, 0, 0) c132176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132176));
	wire w136176;
	repeater #(4, 1'b0, 0, 0) c136176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136176));
	wire w140176;
	repeater #(4, 1'b0, 0, 0) c140176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140176));
	wire w144176;
	repeater #(4, 1'b0, 0, 0) c144176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144176));
	wire w148176;
	repeater #(4, 1'b0, 0, 0) c148176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148176));
	wire w124180;
	repeater #(4, 1'b0, 0, 0) c124180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124180));
	wire w128180;
	repeater #(4, 1'b0, 0, 0) c128180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128180));
	wire w132180;
	repeater #(4, 1'b0, 0, 0) c132180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132180));
	wire w136180;
	repeater #(4, 1'b0, 0, 0) c136180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136180));
	wire w140180;
	repeater #(4, 1'b0, 0, 0) c140180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140180));
	wire w144180;
	repeater #(4, 1'b0, 0, 0) c144180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144180));
	wire w148180;
	repeater #(4, 1'b0, 0, 0) c148180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148180));
	wire w124181;
	repeater #(4, 1'b0, 0, 0) c124181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124181));
	wire w128181;
	repeater #(4, 1'b0, 0, 0) c128181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128181));
	wire w132181;
	repeater #(4, 1'b0, 0, 0) c132181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132181));
	wire w136181;
	repeater #(4, 1'b0, 0, 0) c136181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136181));
	wire w140181;
	repeater #(4, 1'b0, 0, 0) c140181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140181));
	wire w144181;
	repeater #(4, 1'b0, 0, 0) c144181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144181));
	wire w148181;
	repeater #(4, 1'b0, 0, 0) c148181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148181));
	wire w124182;
	repeater #(4, 1'b0, 0, 0) c124182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124182));
	wire w128182;
	repeater #(4, 1'b0, 0, 0) c128182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128182));
	wire w132182;
	repeater #(4, 1'b0, 0, 0) c132182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132182));
	wire w136182;
	repeater #(4, 1'b0, 0, 0) c136182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136182));
	wire w140182;
	repeater #(4, 1'b0, 0, 0) c140182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140182));
	wire w144182;
	repeater #(4, 1'b0, 0, 0) c144182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144182));
	wire w148182;
	repeater #(4, 1'b0, 0, 0) c148182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148182));
	wire w124183;
	repeater #(4, 1'b0, 0, 0) c124183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124183));
	wire w128183;
	repeater #(4, 1'b0, 0, 0) c128183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128183));
	wire w132183;
	repeater #(4, 1'b0, 0, 0) c132183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132183));
	wire w136183;
	repeater #(4, 1'b0, 0, 0) c136183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136183));
	wire w140183;
	repeater #(4, 1'b0, 0, 0) c140183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140183));
	wire w144183;
	repeater #(4, 1'b0, 0, 0) c144183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144183));
	wire w148183;
	repeater #(4, 1'b0, 0, 0) c148183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148183));
	wire w124184;
	repeater #(4, 1'b0, 0, 0) c124184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124184));
	wire w128184;
	repeater #(4, 1'b0, 0, 0) c128184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128184));
	wire w132184;
	repeater #(4, 1'b0, 0, 0) c132184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132184));
	wire w136184;
	repeater #(4, 1'b0, 0, 0) c136184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136184));
	wire w140184;
	repeater #(4, 1'b0, 0, 0) c140184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140184));
	wire w144184;
	repeater #(4, 1'b0, 0, 0) c144184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144184));
	wire w148184;
	repeater #(4, 1'b0, 0, 0) c148184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148184));
	wire w124185;
	repeater #(4, 1'b0, 0, 0) c124185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124185));
	wire w128185;
	repeater #(4, 1'b0, 0, 0) c128185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128185));
	wire w132185;
	repeater #(4, 1'b0, 0, 0) c132185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132185));
	wire w136185;
	repeater #(4, 1'b0, 0, 0) c136185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136185));
	wire w140185;
	repeater #(4, 1'b0, 0, 0) c140185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140185));
	wire w144185;
	repeater #(4, 1'b0, 0, 0) c144185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144185));
	wire w148185;
	repeater #(4, 1'b0, 0, 0) c148185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148185));
	wire w124186;
	repeater #(4, 1'b0, 0, 0) c124186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124186));
	wire w128186;
	repeater #(4, 1'b0, 0, 0) c128186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128186));
	wire w132186;
	repeater #(4, 1'b0, 0, 0) c132186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132186));
	wire w136186;
	repeater #(4, 1'b0, 0, 0) c136186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136186));
	wire w140186;
	repeater #(4, 1'b0, 0, 0) c140186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140186));
	wire w144186;
	repeater #(4, 1'b0, 0, 0) c144186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144186));
	wire w148186;
	repeater #(4, 1'b0, 0, 0) c148186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148186));
	wire w124187;
	repeater #(4, 1'b0, 0, 0) c124187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124187));
	wire w128187;
	repeater #(4, 1'b0, 0, 0) c128187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128187));
	wire w132187;
	repeater #(4, 1'b0, 0, 0) c132187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132187));
	wire w136187;
	repeater #(4, 1'b0, 0, 0) c136187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136187));
	wire w140187;
	repeater #(4, 1'b0, 0, 0) c140187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140187));
	wire w144187;
	repeater #(4, 1'b0, 0, 0) c144187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144187));
	wire w148187;
	repeater #(4, 1'b0, 0, 0) c148187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148187));
	wire w124188;
	repeater #(4, 1'b0, 0, 0) c124188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124188));
	wire w128188;
	repeater #(4, 1'b0, 0, 0) c128188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128188));
	wire w132188;
	repeater #(4, 1'b0, 0, 0) c132188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132188));
	wire w136188;
	repeater #(4, 1'b0, 0, 0) c136188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136188));
	wire w140188;
	repeater #(4, 1'b0, 0, 0) c140188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140188));
	wire w144188;
	repeater #(4, 1'b0, 0, 0) c144188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144188));
	wire w148188;
	repeater #(4, 1'b0, 0, 0) c148188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148188));
	wire w124189;
	repeater #(4, 1'b0, 0, 0) c124189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124189));
	wire w128189;
	repeater #(4, 1'b0, 0, 0) c128189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128189));
	wire w132189;
	repeater #(4, 1'b0, 0, 0) c132189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132189));
	wire w136189;
	repeater #(4, 1'b0, 0, 0) c136189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136189));
	wire w140189;
	repeater #(4, 1'b0, 0, 0) c140189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140189));
	wire w144189;
	repeater #(4, 1'b0, 0, 0) c144189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144189));
	wire w148189;
	repeater #(4, 1'b0, 0, 0) c148189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148189));
	wire w124190;
	repeater #(4, 1'b0, 0, 0) c124190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124190));
	wire w128190;
	repeater #(4, 1'b0, 0, 0) c128190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128190));
	wire w132190;
	repeater #(4, 1'b0, 0, 0) c132190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132190));
	wire w136190;
	repeater #(4, 1'b0, 0, 0) c136190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136190));
	wire w140190;
	repeater #(4, 1'b0, 0, 0) c140190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140190));
	wire w144190;
	repeater #(4, 1'b0, 0, 0) c144190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144190));
	wire w148190;
	repeater #(4, 1'b0, 0, 0) c148190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148190));
	wire w124191;
	repeater #(4, 1'b0, 0, 0) c124191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124191));
	wire w128191;
	repeater #(4, 1'b0, 0, 0) c128191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128191));
	wire w132191;
	repeater #(4, 1'b0, 0, 0) c132191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132191));
	wire w136191;
	repeater #(4, 1'b0, 0, 0) c136191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136191));
	wire w140191;
	repeater #(4, 1'b0, 0, 0) c140191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140191));
	wire w144191;
	repeater #(4, 1'b0, 0, 0) c144191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144191));
	wire w148191;
	repeater #(4, 1'b0, 0, 0) c148191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148191));
	wire w124192;
	repeater #(4, 1'b0, 0, 0) c124192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124192));
	wire w128192;
	repeater #(4, 1'b0, 0, 0) c128192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128192));
	wire w132192;
	repeater #(4, 1'b0, 0, 0) c132192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132192));
	wire w136192;
	repeater #(4, 1'b0, 0, 0) c136192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136192));
	wire w140192;
	repeater #(4, 1'b0, 0, 0) c140192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140192));
	wire w144192;
	repeater #(4, 1'b0, 0, 0) c144192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144192));
	wire w148192;
	repeater #(4, 1'b0, 0, 0) c148192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148192));
	wire w124193;
	repeater #(4, 1'b0, 0, 0) c124193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124193));
	wire w128193;
	repeater #(4, 1'b0, 0, 0) c128193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128193));
	wire w132193;
	repeater #(4, 1'b0, 0, 0) c132193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132193));
	wire w136193;
	repeater #(4, 1'b0, 0, 0) c136193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136193));
	wire w140193;
	repeater #(4, 1'b0, 0, 0) c140193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140193));
	wire w144193;
	repeater #(4, 1'b0, 0, 0) c144193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144193));
	wire w148193;
	repeater #(4, 1'b0, 0, 0) c148193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148193));
	wire w124194;
	repeater #(4, 1'b0, 0, 0) c124194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124194));
	wire w128194;
	repeater #(4, 1'b0, 0, 0) c128194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128194));
	wire w132194;
	repeater #(4, 1'b0, 0, 0) c132194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132194));
	wire w136194;
	repeater #(4, 1'b0, 0, 0) c136194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136194));
	wire w140194;
	repeater #(4, 1'b0, 0, 0) c140194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140194));
	wire w144194;
	repeater #(4, 1'b0, 0, 0) c144194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144194));
	wire w148194;
	repeater #(4, 1'b0, 0, 0) c148194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148194));
	wire w124195;
	repeater #(4, 1'b0, 0, 0) c124195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124195));
	wire w128195;
	repeater #(4, 1'b0, 0, 0) c128195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128195));
	wire w132195;
	repeater #(4, 1'b0, 0, 0) c132195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132195));
	wire w136195;
	repeater #(4, 1'b0, 0, 0) c136195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136195));
	wire w140195;
	repeater #(4, 1'b0, 0, 0) c140195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140195));
	wire w144195;
	repeater #(4, 1'b0, 0, 0) c144195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144195));
	wire w148195;
	repeater #(4, 1'b0, 0, 0) c148195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148195));
	wire w124196;
	repeater #(4, 1'b0, 0, 0) c124196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124196));
	wire w128196;
	repeater #(4, 1'b0, 0, 0) c128196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128196));
	wire w132196;
	repeater #(4, 1'b0, 0, 0) c132196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132196));
	wire w136196;
	repeater #(4, 1'b0, 0, 0) c136196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136196));
	wire w140196;
	repeater #(4, 1'b0, 0, 0) c140196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140196));
	wire w144196;
	repeater #(4, 1'b0, 0, 0) c144196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144196));
	wire w148196;
	repeater #(4, 1'b0, 0, 0) c148196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148196));
	wire w124197;
	repeater #(4, 1'b0, 0, 0) c124197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124197));
	wire w128197;
	repeater #(4, 1'b0, 0, 0) c128197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128197));
	wire w132197;
	repeater #(4, 1'b0, 0, 0) c132197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132197));
	wire w136197;
	repeater #(4, 1'b0, 0, 0) c136197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136197));
	wire w140197;
	repeater #(4, 1'b0, 0, 0) c140197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140197));
	wire w144197;
	repeater #(4, 1'b0, 0, 0) c144197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144197));
	wire w148197;
	repeater #(4, 1'b0, 0, 0) c148197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148197));
	wire w124198;
	repeater #(4, 1'b0, 0, 0) c124198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124198));
	wire w128198;
	repeater #(4, 1'b0, 0, 0) c128198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128198));
	wire w132198;
	repeater #(4, 1'b0, 0, 0) c132198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132198));
	wire w136198;
	repeater #(4, 1'b0, 0, 0) c136198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136198));
	wire w140198;
	repeater #(4, 1'b0, 0, 0) c140198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140198));
	wire w144198;
	repeater #(4, 1'b0, 0, 0) c144198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144198));
	wire w148198;
	repeater #(4, 1'b0, 0, 0) c148198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148198));
	wire w124199;
	repeater #(4, 1'b0, 0, 0) c124199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124199));
	wire w128199;
	repeater #(4, 1'b0, 0, 0) c128199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128199));
	wire w132199;
	repeater #(4, 1'b0, 0, 0) c132199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132199));
	wire w136199;
	repeater #(4, 1'b0, 0, 0) c136199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136199));
	wire w140199;
	repeater #(4, 1'b0, 0, 0) c140199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140199));
	wire w144199;
	repeater #(4, 1'b0, 0, 0) c144199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144199));
	wire w148199;
	repeater #(4, 1'b0, 0, 0) c148199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w148199));
	wire w1241100;
	repeater #(4, 1'b0, 0, 0) c1241100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241100));
	wire w1281100;
	repeater #(4, 1'b0, 0, 0) c1281100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281100));
	wire w1321100;
	repeater #(4, 1'b0, 0, 0) c1321100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321100));
	wire w1361100;
	repeater #(4, 1'b0, 0, 0) c1361100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361100));
	wire w1401100;
	repeater #(4, 1'b0, 0, 0) c1401100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401100));
	wire w1441100;
	repeater #(4, 1'b0, 0, 0) c1441100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441100));
	wire w1481100;
	repeater #(4, 1'b0, 0, 0) c1481100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1481100));
	wire w1241101;
	repeater #(4, 1'b0, 0, 0) c1241101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241101));
	wire w1281101;
	repeater #(4, 1'b0, 0, 0) c1281101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281101));
	wire w1321101;
	repeater #(4, 1'b0, 0, 0) c1321101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321101));
	wire w1361101;
	repeater #(4, 1'b0, 0, 0) c1361101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361101));
	wire w1401101;
	repeater #(4, 1'b0, 0, 0) c1401101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401101));
	wire w1441101;
	repeater #(4, 1'b0, 0, 0) c1441101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441101));
	wire w1481101;
	repeater #(4, 1'b0, 0, 0) c1481101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1481101));
	wire w1201106;
	repeater #(1, 1'b0, 0, 0) c1201106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201106));
	wire w1241106;
	repeater #(1, 1'b0, 0, 0) c1241106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241106));
	wire w1281106;
	repeater #(1, 1'b0, 0, 0) c1281106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281106));
	wire w1321106;
	repeater #(1, 1'b0, 0, 0) c1321106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321106));
	wire w1361106;
	repeater #(1, 1'b0, 0, 0) c1361106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1361106));
	wire w1401106;
	repeater #(1, 1'b0, 0, 0) c1401106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1401106));
	wire w1441106;
	repeater #(1, 1'b0, 0, 0) c1441106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1441106));
	wire w1531121;
	assign outputs[116] = ();
	wire w105022;
	torch #(1'b1) c105022 (.i_clk(tick), .i_in(), .o_out(w105022));
	wire w99034;

	wire w101034;

	wire w100035;
	repeater #(1, 1'b0, 0, 0) c100035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100035));
	wire w65049;
	repeater #(1, 1'b1, 0, 0) c65049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w65049));
	wire w207071;
	repeater #(1, 1'b0, 0, 0) c207071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207071));
	wire w1080155;
	repeater #(1, 1'b0, 0, 0) c1080155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1080155));
	wire w1120155;
	repeater #(1, 1'b0, 0, 0) c1120155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1120155));
	wire w1160155;
	repeater #(1, 1'b0, 0, 0) c1160155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1160155));
	wire w1200155;
	repeater #(1, 1'b0, 0, 0) c1200155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1200155));
	wire w1240155;
	repeater #(1, 1'b0, 0, 0) c1240155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240155));
	wire w1280155;
	repeater #(1, 1'b0, 0, 0) c1280155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1280155));
	wire w1320155;
	repeater #(1, 1'b0, 0, 0) c1320155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1320155));
	wire w1370160;
	repeater #(1, 1'b0, 0, 0) c1370160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370160));
	wire w1390160;

	wire w1400160;
	repeater #(4, 1'b0, 0, 0) c1400160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1400160));
	wire w1390161;
	repeater #(1, 1'b0, 0, 0) c1390161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390161));
	wire w1400162;
	repeater #(4, 1'b0, 0, 0) c1400162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1400162));
	wire w89120;
	repeater #(1, 1'b0, 0, 0) c89120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89120));
	wire w136121;
	repeater #(1, 1'b1, 0, 0) c136121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w136121));
	wire w119122;
	repeater #(1, 1'b1, 0, 0) c119122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119122));
	wire w99125;
	repeater #(1, 1'b0, 0, 0) c99125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99125));
	wire w101125;
	repeater #(1, 1'b0, 0, 0) c101125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101125));
	wire w99126;
	repeater #(2, 1'b0, 0, 0) c99126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99126));
	wire w101126;
	repeater #(2, 1'b0, 0, 0) c101126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101126));
	wire w99127;
	repeater #(2, 1'b0, 0, 0) c99127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99127));
	wire w101127;
	repeater #(2, 1'b0, 0, 0) c101127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101127));
	wire w99128;
	repeater #(2, 1'b0, 0, 0) c99128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99128));
	wire w101128;
	repeater #(2, 1'b0, 0, 0) c101128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101128));
	wire w99129;
	repeater #(2, 1'b0, 0, 0) c99129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99129));
	wire w101129;
	repeater #(2, 1'b0, 0, 0) c101129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w101129));
	wire w108131;
	repeater #(3, 1'b0, 0, 0) c108131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108131));
	wire w112131;
	repeater #(3, 1'b0, 0, 0) c112131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112131));
	wire w116131;
	repeater #(3, 1'b0, 0, 0) c116131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116131));
	wire w120131;
	repeater #(3, 1'b0, 0, 0) c120131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120131));
	wire w124131;
	repeater #(3, 1'b0, 0, 0) c124131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124131));
	wire w128131;
	repeater #(3, 1'b0, 0, 0) c128131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128131));
	wire w132131;
	repeater #(3, 1'b0, 0, 0) c132131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132131));
	wire w107132;
	torch #(1'b0) c107132 (.i_clk(tick), .i_in(), .o_out(w107132));
	wire w111132;
	torch #(1'b0) c111132 (.i_clk(tick), .i_in(), .o_out(w111132));
	wire w115132;
	torch #(1'b0) c115132 (.i_clk(tick), .i_in(), .o_out(w115132));
	wire w119132;
	torch #(1'b0) c119132 (.i_clk(tick), .i_in(), .o_out(w119132));
	wire w123132;
	torch #(1'b0) c123132 (.i_clk(tick), .i_in(), .o_out(w123132));
	wire w127132;
	torch #(1'b0) c127132 (.i_clk(tick), .i_in(), .o_out(w127132));
	wire w131132;
	torch #(1'b0) c131132 (.i_clk(tick), .i_in(), .o_out(w131132));
	wire w103133;
	repeater #(2, 1'b0, 0, 0) c103133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103133));
	wire w103134;
	repeater #(2, 1'b0, 0, 0) c103134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103134));
	wire w103135;
	repeater #(2, 1'b0, 0, 0) c103135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103135));
	wire w108135;
	repeater #(2, 1'b0, 0, 0) c108135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108135));
	wire w112135;
	repeater #(2, 1'b0, 0, 0) c112135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112135));
	wire w116135;
	repeater #(2, 1'b0, 0, 0) c116135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116135));
	wire w120135;
	repeater #(2, 1'b0, 0, 0) c120135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120135));
	wire w124135;
	repeater #(2, 1'b0, 0, 0) c124135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124135));
	wire w128135;
	repeater #(2, 1'b0, 0, 0) c128135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128135));
	wire w132135;
	repeater #(2, 1'b0, 0, 0) c132135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132135));
	wire w103136;
	repeater #(2, 1'b0, 0, 0) c103136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103136));
	wire w108136;
	repeater #(3, 1'b0, 0, 0) c108136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108136));
	wire w112136;
	repeater #(3, 1'b0, 0, 0) c112136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112136));
	wire w116136;
	repeater #(3, 1'b0, 0, 0) c116136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116136));
	wire w120136;
	repeater #(3, 1'b0, 0, 0) c120136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120136));
	wire w124136;
	repeater #(3, 1'b0, 0, 0) c124136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124136));
	wire w128136;
	repeater #(3, 1'b0, 0, 0) c128136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128136));
	wire w132136;
	repeater #(3, 1'b0, 0, 0) c132136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132136));
	wire w103137;
	repeater #(1, 1'b0, 0, 0) c103137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w103137));
	wire w108137;
	repeater #(4, 1'b0, 0, 0) c108137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108137));
	wire w112137;
	repeater #(4, 1'b0, 0, 0) c112137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112137));
	wire w116137;
	repeater #(4, 1'b0, 0, 0) c116137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116137));
	wire w120137;
	repeater #(4, 1'b0, 0, 0) c120137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120137));
	wire w124137;
	repeater #(4, 1'b0, 0, 0) c124137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124137));
	wire w128137;
	repeater #(4, 1'b0, 0, 0) c128137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128137));
	wire w132137;
	repeater #(4, 1'b0, 0, 0) c132137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132137));
	wire w108138;
	repeater #(4, 1'b0, 0, 0) c108138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108138));
	wire w112138;
	repeater #(4, 1'b0, 0, 0) c112138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112138));
	wire w116138;
	repeater #(4, 1'b0, 0, 0) c116138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116138));
	wire w120138;
	repeater #(4, 1'b0, 0, 0) c120138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120138));
	wire w124138;
	repeater #(4, 1'b0, 0, 0) c124138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124138));
	wire w128138;
	repeater #(4, 1'b0, 0, 0) c128138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128138));
	wire w132138;
	repeater #(4, 1'b0, 0, 0) c132138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132138));
	wire w108139;
	repeater #(4, 1'b0, 0, 0) c108139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108139));
	wire w112139;
	repeater #(4, 1'b0, 0, 0) c112139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112139));
	wire w116139;
	repeater #(4, 1'b0, 0, 0) c116139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116139));
	wire w120139;
	repeater #(4, 1'b0, 0, 0) c120139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120139));
	wire w124139;
	repeater #(4, 1'b0, 0, 0) c124139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124139));
	wire w128139;
	repeater #(4, 1'b0, 0, 0) c128139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128139));
	wire w132139;
	repeater #(4, 1'b0, 0, 0) c132139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132139));
	wire w108140;
	repeater #(4, 1'b0, 0, 0) c108140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108140));
	wire w112140;
	repeater #(4, 1'b0, 0, 0) c112140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112140));
	wire w116140;
	repeater #(4, 1'b0, 0, 0) c116140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116140));
	wire w120140;
	repeater #(4, 1'b0, 0, 0) c120140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120140));
	wire w124140;
	repeater #(4, 1'b0, 0, 0) c124140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124140));
	wire w128140;
	repeater #(4, 1'b0, 0, 0) c128140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128140));
	wire w132140;
	repeater #(4, 1'b0, 0, 0) c132140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132140));
	wire w108141;
	repeater #(4, 1'b0, 0, 0) c108141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108141));
	wire w112141;
	repeater #(4, 1'b0, 0, 0) c112141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112141));
	wire w116141;
	repeater #(4, 1'b0, 0, 0) c116141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116141));
	wire w120141;
	repeater #(4, 1'b0, 0, 0) c120141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120141));
	wire w124141;
	repeater #(4, 1'b0, 0, 0) c124141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124141));
	wire w128141;
	repeater #(4, 1'b0, 0, 0) c128141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128141));
	wire w132141;
	repeater #(4, 1'b0, 0, 0) c132141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132141));
	wire w108142;
	repeater #(4, 1'b0, 0, 0) c108142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108142));
	wire w112142;
	repeater #(4, 1'b0, 0, 0) c112142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112142));
	wire w116142;
	repeater #(4, 1'b0, 0, 0) c116142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116142));
	wire w120142;
	repeater #(4, 1'b0, 0, 0) c120142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120142));
	wire w124142;
	repeater #(4, 1'b0, 0, 0) c124142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124142));
	wire w128142;
	repeater #(4, 1'b0, 0, 0) c128142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128142));
	wire w132142;
	repeater #(4, 1'b0, 0, 0) c132142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132142));
	wire w108143;
	repeater #(4, 1'b0, 0, 0) c108143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108143));
	wire w112143;
	repeater #(4, 1'b0, 0, 0) c112143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112143));
	wire w116143;
	repeater #(4, 1'b0, 0, 0) c116143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116143));
	wire w120143;
	repeater #(4, 1'b0, 0, 0) c120143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120143));
	wire w124143;
	repeater #(4, 1'b0, 0, 0) c124143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124143));
	wire w128143;
	repeater #(4, 1'b0, 0, 0) c128143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128143));
	wire w132143;
	repeater #(4, 1'b0, 0, 0) c132143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132143));
	wire w108144;
	repeater #(4, 1'b0, 0, 0) c108144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108144));
	wire w112144;
	repeater #(4, 1'b0, 0, 0) c112144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112144));
	wire w116144;
	repeater #(4, 1'b0, 0, 0) c116144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116144));
	wire w120144;
	repeater #(4, 1'b0, 0, 0) c120144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120144));
	wire w124144;
	repeater #(4, 1'b0, 0, 0) c124144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124144));
	wire w128144;
	repeater #(4, 1'b0, 0, 0) c128144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128144));
	wire w132144;
	repeater #(4, 1'b0, 0, 0) c132144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132144));
	wire w108145;
	repeater #(4, 1'b0, 0, 0) c108145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108145));
	wire w112145;
	repeater #(4, 1'b0, 0, 0) c112145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112145));
	wire w116145;
	repeater #(4, 1'b0, 0, 0) c116145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116145));
	wire w120145;
	repeater #(4, 1'b0, 0, 0) c120145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120145));
	wire w124145;
	repeater #(4, 1'b0, 0, 0) c124145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124145));
	wire w128145;
	repeater #(4, 1'b0, 0, 0) c128145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128145));
	wire w132145;
	repeater #(4, 1'b0, 0, 0) c132145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132145));
	wire w108146;
	repeater #(4, 1'b0, 0, 0) c108146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108146));
	wire w112146;
	repeater #(4, 1'b0, 0, 0) c112146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112146));
	wire w116146;
	repeater #(4, 1'b0, 0, 0) c116146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116146));
	wire w120146;
	repeater #(4, 1'b0, 0, 0) c120146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120146));
	wire w124146;
	repeater #(4, 1'b0, 0, 0) c124146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124146));
	wire w128146;
	repeater #(4, 1'b0, 0, 0) c128146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128146));
	wire w132146;
	repeater #(4, 1'b0, 0, 0) c132146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132146));
	wire w108147;
	repeater #(4, 1'b0, 0, 0) c108147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108147));
	wire w112147;
	repeater #(4, 1'b0, 0, 0) c112147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112147));
	wire w116147;
	repeater #(4, 1'b0, 0, 0) c116147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116147));
	wire w120147;
	repeater #(4, 1'b0, 0, 0) c120147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120147));
	wire w124147;
	repeater #(4, 1'b0, 0, 0) c124147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124147));
	wire w128147;
	repeater #(4, 1'b0, 0, 0) c128147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128147));
	wire w132147;
	repeater #(4, 1'b0, 0, 0) c132147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132147));
	wire w66148;

	wire w108148;
	repeater #(4, 1'b0, 0, 0) c108148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108148));
	wire w112148;
	repeater #(4, 1'b0, 0, 0) c112148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112148));
	wire w116148;
	repeater #(4, 1'b0, 0, 0) c116148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116148));
	wire w120148;
	repeater #(4, 1'b0, 0, 0) c120148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120148));
	wire w124148;
	repeater #(4, 1'b0, 0, 0) c124148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124148));
	wire w128148;
	repeater #(4, 1'b0, 0, 0) c128148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128148));
	wire w132148;
	repeater #(4, 1'b0, 0, 0) c132148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132148));
	wire w108149;
	repeater #(2, 1'b0, 0, 0) c108149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108149));
	wire w112149;
	repeater #(2, 1'b0, 0, 0) c112149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112149));
	wire w116149;
	repeater #(2, 1'b0, 0, 0) c116149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116149));
	wire w120149;
	repeater #(2, 1'b0, 0, 0) c120149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120149));
	wire w124149;
	repeater #(2, 1'b0, 0, 0) c124149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124149));
	wire w128149;
	repeater #(2, 1'b0, 0, 0) c128149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128149));
	wire w132149;
	repeater #(2, 1'b0, 0, 0) c132149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132149));
	wire w133153;
	repeater #(2, 1'b1, 0, 0) c133153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133153));
	wire w107154;
	repeater #(2, 1'b1, 0, 0) c107154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107154));
	wire w108154;
	repeater #(1, 1'b0, 0, 0) c108154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108154));
	wire w111154;
	repeater #(2, 1'b1, 0, 0) c111154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111154));
	wire w112154;
	repeater #(1, 1'b0, 0, 0) c112154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112154));
	wire w115154;
	repeater #(2, 1'b1, 0, 0) c115154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115154));
	wire w116154;
	repeater #(1, 1'b0, 0, 0) c116154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116154));
	wire w119154;
	repeater #(2, 1'b1, 0, 0) c119154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119154));
	wire w120154;
	repeater #(1, 1'b0, 0, 0) c120154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120154));
	wire w123154;
	repeater #(2, 1'b1, 0, 0) c123154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123154));
	wire w124154;
	repeater #(1, 1'b0, 0, 0) c124154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124154));
	wire w127154;
	repeater #(2, 1'b1, 0, 0) c127154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127154));
	wire w128154;
	repeater #(1, 1'b0, 0, 0) c128154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128154));
	wire w131154;
	repeater #(2, 1'b1, 0, 0) c131154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131154));
	wire w132154;
	repeater #(1, 1'b0, 0, 0) c132154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132154));
	wire w107155;
	torch #(1'b0) c107155 (.i_clk(tick), .i_in(), .o_out(w107155));
	wire w111155;
	torch #(1'b0) c111155 (.i_clk(tick), .i_in(), .o_out(w111155));
	wire w115155;
	torch #(1'b0) c115155 (.i_clk(tick), .i_in(), .o_out(w115155));
	wire w119155;
	torch #(1'b0) c119155 (.i_clk(tick), .i_in(), .o_out(w119155));
	wire w123155;
	torch #(1'b0) c123155 (.i_clk(tick), .i_in(), .o_out(w123155));
	wire w127155;
	torch #(1'b0) c127155 (.i_clk(tick), .i_in(), .o_out(w127155));
	wire w131155;
	torch #(1'b0) c131155 (.i_clk(tick), .i_in(), .o_out(w131155));
	wire w108156;
	repeater #(4, 1'b0, 0, 0) c108156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108156));
	wire w112156;
	repeater #(4, 1'b0, 0, 0) c112156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112156));
	wire w116156;
	repeater #(4, 1'b0, 0, 0) c116156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116156));
	wire w120156;
	repeater #(4, 1'b0, 0, 0) c120156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120156));
	wire w124156;
	repeater #(4, 1'b0, 0, 0) c124156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124156));
	wire w128156;
	repeater #(4, 1'b0, 0, 0) c128156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128156));
	wire w132156;
	repeater #(4, 1'b0, 0, 0) c132156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132156));
	wire w108157;
	repeater #(4, 1'b0, 0, 0) c108157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108157));
	wire w112157;
	repeater #(4, 1'b0, 0, 0) c112157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112157));
	wire w116157;
	repeater #(4, 1'b0, 0, 0) c116157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116157));
	wire w120157;
	repeater #(4, 1'b0, 0, 0) c120157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120157));
	wire w124157;
	repeater #(4, 1'b0, 0, 0) c124157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124157));
	wire w128157;
	repeater #(4, 1'b0, 0, 0) c128157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128157));
	wire w132157;
	repeater #(4, 1'b0, 0, 0) c132157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132157));
	wire w138157;
	repeater #(1, 1'b1, 0, 0) c138157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138157));
	wire w140157;
	repeater #(1, 1'b1, 0, 0) c140157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140157));
	wire w142157;
	repeater #(1, 1'b1, 0, 0) c142157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142157));
	wire w108158;
	repeater #(4, 1'b0, 0, 0) c108158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108158));
	wire w112158;
	repeater #(4, 1'b0, 0, 0) c112158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112158));
	wire w116158;
	repeater #(4, 1'b0, 0, 0) c116158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116158));
	wire w120158;
	repeater #(4, 1'b0, 0, 0) c120158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120158));
	wire w124158;
	repeater #(4, 1'b0, 0, 0) c124158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124158));
	wire w128158;
	repeater #(4, 1'b0, 0, 0) c128158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128158));
	wire w132158;
	repeater #(4, 1'b0, 0, 0) c132158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132158));
	wire w108159;
	repeater #(4, 1'b0, 0, 0) c108159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108159));
	wire w112159;
	repeater #(4, 1'b0, 0, 0) c112159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112159));
	wire w116159;
	repeater #(4, 1'b0, 0, 0) c116159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116159));
	wire w120159;
	repeater #(4, 1'b0, 0, 0) c120159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120159));
	wire w124159;
	repeater #(4, 1'b0, 0, 0) c124159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124159));
	wire w128159;
	repeater #(4, 1'b0, 0, 0) c128159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128159));
	wire w132159;
	repeater #(4, 1'b0, 0, 0) c132159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132159));
	wire w108160;
	repeater #(4, 1'b0, 0, 0) c108160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108160));
	wire w112160;
	repeater #(4, 1'b0, 0, 0) c112160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112160));
	wire w116160;
	repeater #(4, 1'b0, 0, 0) c116160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116160));
	wire w120160;
	repeater #(4, 1'b0, 0, 0) c120160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120160));
	wire w124160;
	repeater #(4, 1'b0, 0, 0) c124160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124160));
	wire w128160;
	repeater #(4, 1'b0, 0, 0) c128160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128160));
	wire w132160;
	repeater #(4, 1'b0, 0, 0) c132160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132160));
	wire w108161;
	repeater #(4, 1'b0, 0, 0) c108161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108161));
	wire w112161;
	repeater #(4, 1'b0, 0, 0) c112161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112161));
	wire w116161;
	repeater #(4, 1'b0, 0, 0) c116161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116161));
	wire w120161;
	repeater #(4, 1'b0, 0, 0) c120161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120161));
	wire w124161;
	repeater #(4, 1'b0, 0, 0) c124161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124161));
	wire w128161;
	repeater #(4, 1'b0, 0, 0) c128161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128161));
	wire w132161;
	repeater #(4, 1'b0, 0, 0) c132161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132161));
	wire w108162;
	repeater #(4, 1'b0, 0, 0) c108162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108162));
	wire w112162;
	repeater #(4, 1'b0, 0, 0) c112162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112162));
	wire w116162;
	repeater #(4, 1'b0, 0, 0) c116162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116162));
	wire w120162;
	repeater #(4, 1'b0, 0, 0) c120162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120162));
	wire w124162;
	repeater #(4, 1'b0, 0, 0) c124162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124162));
	wire w128162;
	repeater #(4, 1'b0, 0, 0) c128162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128162));
	wire w132162;
	repeater #(4, 1'b0, 0, 0) c132162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132162));
	wire w108163;
	repeater #(4, 1'b0, 0, 0) c108163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108163));
	wire w112163;
	repeater #(4, 1'b0, 0, 0) c112163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112163));
	wire w116163;
	repeater #(4, 1'b0, 0, 0) c116163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116163));
	wire w120163;
	repeater #(4, 1'b0, 0, 0) c120163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120163));
	wire w124163;
	repeater #(4, 1'b0, 0, 0) c124163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124163));
	wire w128163;
	repeater #(4, 1'b0, 0, 0) c128163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128163));
	wire w132163;
	repeater #(4, 1'b0, 0, 0) c132163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132163));
	wire w108164;
	repeater #(4, 1'b0, 0, 0) c108164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108164));
	wire w112164;
	repeater #(4, 1'b0, 0, 0) c112164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112164));
	wire w116164;
	repeater #(4, 1'b0, 0, 0) c116164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116164));
	wire w120164;
	repeater #(4, 1'b0, 0, 0) c120164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120164));
	wire w124164;
	repeater #(4, 1'b0, 0, 0) c124164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124164));
	wire w128164;
	repeater #(4, 1'b0, 0, 0) c128164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128164));
	wire w132164;
	repeater #(4, 1'b0, 0, 0) c132164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132164));
	wire w108165;
	repeater #(4, 1'b0, 0, 0) c108165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108165));
	wire w112165;
	repeater #(4, 1'b0, 0, 0) c112165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112165));
	wire w116165;
	repeater #(4, 1'b0, 0, 0) c116165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116165));
	wire w120165;
	repeater #(4, 1'b0, 0, 0) c120165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120165));
	wire w124165;
	repeater #(4, 1'b0, 0, 0) c124165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124165));
	wire w128165;
	repeater #(4, 1'b0, 0, 0) c128165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128165));
	wire w132165;
	repeater #(4, 1'b0, 0, 0) c132165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132165));
	wire w108166;
	repeater #(4, 1'b0, 0, 0) c108166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108166));
	wire w112166;
	repeater #(4, 1'b0, 0, 0) c112166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112166));
	wire w116166;
	repeater #(4, 1'b0, 0, 0) c116166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116166));
	wire w120166;
	repeater #(4, 1'b0, 0, 0) c120166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120166));
	wire w124166;
	repeater #(4, 1'b0, 0, 0) c124166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124166));
	wire w128166;
	repeater #(4, 1'b0, 0, 0) c128166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128166));
	wire w132166;
	repeater #(4, 1'b0, 0, 0) c132166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132166));
	wire w108167;
	repeater #(4, 1'b0, 0, 0) c108167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108167));
	wire w112167;
	repeater #(4, 1'b0, 0, 0) c112167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112167));
	wire w116167;
	repeater #(4, 1'b0, 0, 0) c116167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116167));
	wire w120167;
	repeater #(4, 1'b0, 0, 0) c120167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120167));
	wire w124167;
	repeater #(4, 1'b0, 0, 0) c124167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124167));
	wire w128167;
	repeater #(4, 1'b0, 0, 0) c128167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128167));
	wire w132167;
	repeater #(4, 1'b0, 0, 0) c132167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132167));
	wire w108168;
	repeater #(4, 1'b0, 0, 0) c108168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108168));
	wire w112168;
	repeater #(4, 1'b0, 0, 0) c112168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112168));
	wire w116168;
	repeater #(4, 1'b0, 0, 0) c116168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116168));
	wire w120168;
	repeater #(4, 1'b0, 0, 0) c120168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120168));
	wire w124168;
	repeater #(4, 1'b0, 0, 0) c124168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124168));
	wire w128168;
	repeater #(4, 1'b0, 0, 0) c128168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128168));
	wire w132168;
	repeater #(4, 1'b0, 0, 0) c132168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132168));
	wire w108169;
	repeater #(4, 1'b0, 0, 0) c108169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108169));
	wire w112169;
	repeater #(4, 1'b0, 0, 0) c112169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112169));
	wire w116169;
	repeater #(4, 1'b0, 0, 0) c116169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116169));
	wire w120169;
	repeater #(4, 1'b0, 0, 0) c120169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120169));
	wire w124169;
	repeater #(4, 1'b0, 0, 0) c124169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124169));
	wire w128169;
	repeater #(4, 1'b0, 0, 0) c128169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128169));
	wire w132169;
	repeater #(4, 1'b0, 0, 0) c132169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132169));
	wire w108170;
	repeater #(4, 1'b0, 0, 0) c108170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108170));
	wire w112170;
	repeater #(4, 1'b0, 0, 0) c112170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112170));
	wire w116170;
	repeater #(4, 1'b0, 0, 0) c116170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116170));
	wire w120170;
	repeater #(4, 1'b0, 0, 0) c120170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120170));
	wire w124170;
	repeater #(4, 1'b0, 0, 0) c124170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124170));
	wire w128170;
	repeater #(4, 1'b0, 0, 0) c128170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128170));
	wire w132170;
	repeater #(4, 1'b0, 0, 0) c132170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132170));
	wire w108171;
	repeater #(4, 1'b0, 0, 0) c108171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108171));
	wire w112171;
	repeater #(4, 1'b0, 0, 0) c112171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112171));
	wire w116171;
	repeater #(4, 1'b0, 0, 0) c116171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116171));
	wire w120171;
	repeater #(4, 1'b0, 0, 0) c120171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120171));
	wire w124171;
	repeater #(4, 1'b0, 0, 0) c124171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124171));
	wire w128171;
	repeater #(4, 1'b0, 0, 0) c128171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128171));
	wire w132171;
	repeater #(4, 1'b0, 0, 0) c132171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132171));
	wire w108172;
	repeater #(4, 1'b0, 0, 0) c108172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108172));
	wire w112172;
	repeater #(4, 1'b0, 0, 0) c112172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112172));
	wire w116172;
	repeater #(4, 1'b0, 0, 0) c116172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116172));
	wire w120172;
	repeater #(4, 1'b0, 0, 0) c120172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120172));
	wire w124172;
	repeater #(4, 1'b0, 0, 0) c124172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124172));
	wire w128172;
	repeater #(4, 1'b0, 0, 0) c128172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128172));
	wire w132172;
	repeater #(4, 1'b0, 0, 0) c132172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132172));
	wire w108173;
	repeater #(4, 1'b0, 0, 0) c108173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108173));
	wire w112173;
	repeater #(4, 1'b0, 0, 0) c112173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112173));
	wire w116173;
	repeater #(4, 1'b0, 0, 0) c116173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116173));
	wire w120173;
	repeater #(4, 1'b0, 0, 0) c120173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120173));
	wire w124173;
	repeater #(4, 1'b0, 0, 0) c124173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124173));
	wire w128173;
	repeater #(4, 1'b0, 0, 0) c128173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128173));
	wire w132173;
	repeater #(4, 1'b0, 0, 0) c132173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132173));
	wire w107178;
	repeater #(3, 1'b1, 0, 0) c107178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w107178));
	wire w108178;
	repeater #(1, 1'b0, 0, 0) c108178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108178));
	wire w111178;
	repeater #(3, 1'b1, 0, 0) c111178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w111178));
	wire w112178;
	repeater #(1, 1'b0, 0, 0) c112178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112178));
	wire w115178;
	repeater #(3, 1'b1, 0, 0) c115178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w115178));
	wire w116178;
	repeater #(1, 1'b0, 0, 0) c116178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116178));
	wire w119178;
	repeater #(3, 1'b1, 0, 0) c119178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w119178));
	wire w120178;
	repeater #(1, 1'b0, 0, 0) c120178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120178));
	wire w123178;
	repeater #(3, 1'b1, 0, 0) c123178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123178));
	wire w124178;
	repeater #(1, 1'b0, 0, 0) c124178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124178));
	wire w127178;
	repeater #(3, 1'b1, 0, 0) c127178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127178));
	wire w128178;
	repeater #(1, 1'b0, 0, 0) c128178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128178));
	wire w131178;
	repeater #(3, 1'b1, 0, 0) c131178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w131178));
	wire w132178;
	repeater #(1, 1'b0, 0, 0) c132178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132178));
	wire w107179;
	torch #(1'b0) c107179 (.i_clk(tick), .i_in(), .o_out(w107179));
	wire w111179;
	torch #(1'b0) c111179 (.i_clk(tick), .i_in(), .o_out(w111179));
	wire w115179;
	torch #(1'b0) c115179 (.i_clk(tick), .i_in(), .o_out(w115179));
	wire w119179;
	torch #(1'b0) c119179 (.i_clk(tick), .i_in(), .o_out(w119179));
	wire w123179;
	torch #(1'b0) c123179 (.i_clk(tick), .i_in(), .o_out(w123179));
	wire w127179;
	torch #(1'b0) c127179 (.i_clk(tick), .i_in(), .o_out(w127179));
	wire w131179;
	torch #(1'b0) c131179 (.i_clk(tick), .i_in(), .o_out(w131179));
	wire w108180;
	repeater #(4, 1'b0, 0, 0) c108180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108180));
	wire w112180;
	repeater #(4, 1'b0, 0, 0) c112180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112180));
	wire w116180;
	repeater #(4, 1'b0, 0, 0) c116180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116180));
	wire w120180;
	repeater #(4, 1'b0, 0, 0) c120180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120180));
	wire w124180;
	repeater #(4, 1'b0, 0, 0) c124180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124180));
	wire w128180;
	repeater #(4, 1'b0, 0, 0) c128180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128180));
	wire w132180;
	repeater #(4, 1'b0, 0, 0) c132180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132180));
	wire w108181;
	repeater #(4, 1'b0, 0, 0) c108181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108181));
	wire w112181;
	repeater #(4, 1'b0, 0, 0) c112181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112181));
	wire w116181;
	repeater #(4, 1'b0, 0, 0) c116181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116181));
	wire w120181;
	repeater #(4, 1'b0, 0, 0) c120181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120181));
	wire w124181;
	repeater #(2, 1'b0, 0, 0) c124181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124181));
	wire w128181;
	repeater #(4, 1'b0, 0, 0) c128181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128181));
	wire w132181;
	repeater #(4, 1'b0, 0, 0) c132181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132181));
	wire w108182;
	repeater #(4, 1'b0, 0, 0) c108182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108182));
	wire w112182;
	repeater #(4, 1'b0, 0, 0) c112182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112182));
	wire w116182;
	repeater #(4, 1'b0, 0, 0) c116182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116182));
	wire w120182;
	repeater #(4, 1'b0, 0, 0) c120182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120182));
	wire w124182;
	repeater #(4, 1'b0, 0, 0) c124182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124182));
	wire w128182;
	repeater #(4, 1'b0, 0, 0) c128182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128182));
	wire w132182;
	repeater #(4, 1'b0, 0, 0) c132182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132182));
	wire w108183;
	repeater #(4, 1'b0, 0, 0) c108183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108183));
	wire w112183;
	repeater #(4, 1'b0, 0, 0) c112183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112183));
	wire w116183;
	repeater #(4, 1'b0, 0, 0) c116183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116183));
	wire w120183;
	repeater #(4, 1'b0, 0, 0) c120183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120183));
	wire w124183;
	repeater #(4, 1'b0, 0, 0) c124183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124183));
	wire w128183;
	repeater #(4, 1'b0, 0, 0) c128183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128183));
	wire w132183;
	repeater #(4, 1'b0, 0, 0) c132183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132183));
	wire w108184;
	repeater #(4, 1'b0, 0, 0) c108184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108184));
	wire w112184;
	repeater #(4, 1'b0, 0, 0) c112184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112184));
	wire w116184;
	repeater #(4, 1'b0, 0, 0) c116184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116184));
	wire w120184;
	repeater #(4, 1'b0, 0, 0) c120184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120184));
	wire w124184;
	repeater #(4, 1'b0, 0, 0) c124184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124184));
	wire w128184;
	repeater #(4, 1'b0, 0, 0) c128184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128184));
	wire w132184;
	repeater #(4, 1'b0, 0, 0) c132184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132184));
	wire w108185;
	repeater #(4, 1'b0, 0, 0) c108185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108185));
	wire w112185;
	repeater #(4, 1'b0, 0, 0) c112185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112185));
	wire w116185;
	repeater #(4, 1'b0, 0, 0) c116185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116185));
	wire w120185;
	repeater #(4, 1'b0, 0, 0) c120185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120185));
	wire w124185;
	repeater #(4, 1'b0, 0, 0) c124185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124185));
	wire w128185;
	repeater #(4, 1'b0, 0, 0) c128185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128185));
	wire w132185;
	repeater #(4, 1'b0, 0, 0) c132185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132185));
	wire w108186;
	repeater #(4, 1'b0, 0, 0) c108186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108186));
	wire w112186;
	repeater #(4, 1'b0, 0, 0) c112186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112186));
	wire w116186;
	repeater #(4, 1'b0, 0, 0) c116186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116186));
	wire w120186;
	repeater #(4, 1'b0, 0, 0) c120186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120186));
	wire w124186;
	repeater #(4, 1'b0, 0, 0) c124186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124186));
	wire w128186;
	repeater #(4, 1'b0, 0, 0) c128186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128186));
	wire w132186;
	repeater #(4, 1'b0, 0, 0) c132186 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132186));
	wire w108187;
	repeater #(4, 1'b0, 0, 0) c108187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108187));
	wire w112187;
	repeater #(4, 1'b0, 0, 0) c112187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112187));
	wire w116187;
	repeater #(4, 1'b0, 0, 0) c116187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116187));
	wire w120187;
	repeater #(4, 1'b0, 0, 0) c120187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120187));
	wire w124187;
	repeater #(4, 1'b0, 0, 0) c124187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124187));
	wire w128187;
	repeater #(4, 1'b0, 0, 0) c128187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128187));
	wire w132187;
	repeater #(4, 1'b0, 0, 0) c132187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132187));
	wire w108188;
	repeater #(4, 1'b0, 0, 0) c108188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108188));
	wire w112188;
	repeater #(4, 1'b0, 0, 0) c112188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112188));
	wire w116188;
	repeater #(4, 1'b0, 0, 0) c116188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116188));
	wire w120188;
	repeater #(4, 1'b0, 0, 0) c120188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120188));
	wire w124188;
	repeater #(4, 1'b0, 0, 0) c124188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124188));
	wire w128188;
	repeater #(4, 1'b0, 0, 0) c128188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128188));
	wire w132188;
	repeater #(4, 1'b0, 0, 0) c132188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132188));
	wire w108189;
	repeater #(4, 1'b0, 0, 0) c108189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108189));
	wire w112189;
	repeater #(4, 1'b0, 0, 0) c112189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112189));
	wire w116189;
	repeater #(4, 1'b0, 0, 0) c116189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116189));
	wire w120189;
	repeater #(4, 1'b0, 0, 0) c120189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120189));
	wire w124189;
	repeater #(4, 1'b0, 0, 0) c124189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124189));
	wire w128189;
	repeater #(4, 1'b0, 0, 0) c128189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128189));
	wire w132189;
	repeater #(4, 1'b0, 0, 0) c132189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132189));
	wire w108190;
	repeater #(4, 1'b0, 0, 0) c108190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108190));
	wire w112190;
	repeater #(4, 1'b0, 0, 0) c112190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112190));
	wire w116190;
	repeater #(4, 1'b0, 0, 0) c116190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116190));
	wire w120190;
	repeater #(4, 1'b0, 0, 0) c120190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120190));
	wire w124190;
	repeater #(4, 1'b0, 0, 0) c124190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124190));
	wire w128190;
	repeater #(4, 1'b0, 0, 0) c128190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128190));
	wire w132190;
	repeater #(4, 1'b0, 0, 0) c132190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132190));
	wire w108191;
	repeater #(4, 1'b0, 0, 0) c108191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108191));
	wire w112191;
	repeater #(4, 1'b0, 0, 0) c112191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112191));
	wire w116191;
	repeater #(4, 1'b0, 0, 0) c116191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116191));
	wire w120191;
	repeater #(4, 1'b0, 0, 0) c120191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120191));
	wire w124191;
	repeater #(4, 1'b0, 0, 0) c124191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124191));
	wire w128191;
	repeater #(4, 1'b0, 0, 0) c128191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128191));
	wire w132191;
	repeater #(4, 1'b0, 0, 0) c132191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132191));
	wire w108192;
	repeater #(4, 1'b0, 0, 0) c108192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108192));
	wire w112192;
	repeater #(4, 1'b0, 0, 0) c112192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112192));
	wire w116192;
	repeater #(4, 1'b0, 0, 0) c116192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116192));
	wire w120192;
	repeater #(4, 1'b0, 0, 0) c120192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120192));
	wire w124192;
	repeater #(4, 1'b0, 0, 0) c124192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124192));
	wire w128192;
	repeater #(4, 1'b0, 0, 0) c128192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128192));
	wire w132192;
	repeater #(4, 1'b0, 0, 0) c132192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132192));
	wire w108193;
	repeater #(4, 1'b0, 0, 0) c108193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108193));
	wire w112193;
	repeater #(4, 1'b0, 0, 0) c112193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112193));
	wire w116193;
	repeater #(4, 1'b0, 0, 0) c116193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116193));
	wire w120193;
	repeater #(4, 1'b0, 0, 0) c120193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120193));
	wire w124193;
	repeater #(4, 1'b0, 0, 0) c124193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124193));
	wire w128193;
	repeater #(4, 1'b0, 0, 0) c128193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128193));
	wire w132193;
	repeater #(4, 1'b0, 0, 0) c132193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132193));
	wire w108194;
	repeater #(4, 1'b0, 0, 0) c108194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108194));
	wire w112194;
	repeater #(4, 1'b0, 0, 0) c112194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112194));
	wire w116194;
	repeater #(4, 1'b0, 0, 0) c116194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116194));
	wire w120194;
	repeater #(4, 1'b0, 0, 0) c120194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120194));
	wire w124194;
	repeater #(4, 1'b0, 0, 0) c124194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124194));
	wire w128194;
	repeater #(4, 1'b0, 0, 0) c128194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128194));
	wire w132194;
	repeater #(4, 1'b0, 0, 0) c132194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132194));
	wire w108195;
	repeater #(4, 1'b0, 0, 0) c108195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108195));
	wire w112195;
	repeater #(4, 1'b0, 0, 0) c112195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112195));
	wire w116195;
	repeater #(4, 1'b0, 0, 0) c116195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116195));
	wire w120195;
	repeater #(4, 1'b0, 0, 0) c120195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120195));
	wire w124195;
	repeater #(4, 1'b0, 0, 0) c124195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124195));
	wire w128195;
	repeater #(4, 1'b0, 0, 0) c128195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128195));
	wire w132195;
	repeater #(4, 1'b0, 0, 0) c132195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132195));
	wire w108196;
	repeater #(4, 1'b0, 0, 0) c108196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108196));
	wire w112196;
	repeater #(4, 1'b0, 0, 0) c112196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w112196));
	wire w116196;
	repeater #(4, 1'b0, 0, 0) c116196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116196));
	wire w120196;
	repeater #(4, 1'b0, 0, 0) c120196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120196));
	wire w124196;
	repeater #(4, 1'b0, 0, 0) c124196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124196));
	wire w128196;
	repeater #(4, 1'b0, 0, 0) c128196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w128196));
	wire w132196;
	repeater #(4, 1'b0, 0, 0) c132196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132196));
	wire w1071102;
	repeater #(3, 1'b1, 0, 0) c1071102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1071102));
	wire w1081102;
	repeater #(1, 1'b0, 0, 0) c1081102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081102));
	wire w1111102;
	repeater #(3, 1'b1, 0, 0) c1111102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1111102));
	wire w1121102;
	repeater #(1, 1'b0, 0, 0) c1121102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121102));
	wire w1151102;
	repeater #(3, 1'b1, 0, 0) c1151102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1151102));
	wire w1161102;
	repeater #(1, 1'b0, 0, 0) c1161102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161102));
	wire w1191102;
	repeater #(3, 1'b1, 0, 0) c1191102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1191102));
	wire w1201102;
	repeater #(1, 1'b0, 0, 0) c1201102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201102));
	wire w1231102;
	repeater #(3, 1'b1, 0, 0) c1231102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1231102));
	wire w1241102;
	repeater #(1, 1'b0, 0, 0) c1241102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241102));
	wire w1271102;
	repeater #(3, 1'b1, 0, 0) c1271102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271102));
	wire w1281102;
	repeater #(1, 1'b0, 0, 0) c1281102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281102));
	wire w1311102;
	repeater #(3, 1'b1, 0, 0) c1311102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1311102));
	wire w1321102;
	repeater #(1, 1'b0, 0, 0) c1321102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321102));
	wire w1071103;
	torch #(1'b0) c1071103 (.i_clk(tick), .i_in(), .o_out(w1071103));
	wire w1111103;
	torch #(1'b0) c1111103 (.i_clk(tick), .i_in(), .o_out(w1111103));
	wire w1151103;
	torch #(1'b0) c1151103 (.i_clk(tick), .i_in(), .o_out(w1151103));
	wire w1191103;
	torch #(1'b0) c1191103 (.i_clk(tick), .i_in(), .o_out(w1191103));
	wire w1231103;
	torch #(1'b0) c1231103 (.i_clk(tick), .i_in(), .o_out(w1231103));
	wire w1271103;
	torch #(1'b0) c1271103 (.i_clk(tick), .i_in(), .o_out(w1271103));
	wire w1311103;
	torch #(1'b0) c1311103 (.i_clk(tick), .i_in(), .o_out(w1311103));
	wire w1081104;
	repeater #(4, 1'b0, 0, 0) c1081104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081104));
	wire w1121104;
	repeater #(4, 1'b0, 0, 0) c1121104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121104));
	wire w1161104;
	repeater #(4, 1'b0, 0, 0) c1161104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161104));
	wire w1201104;
	repeater #(4, 1'b0, 0, 0) c1201104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201104));
	wire w1241104;
	repeater #(4, 1'b0, 0, 0) c1241104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241104));
	wire w1281104;
	repeater #(4, 1'b0, 0, 0) c1281104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281104));
	wire w1321104;
	repeater #(4, 1'b0, 0, 0) c1321104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321104));
	wire w1081105;
	repeater #(4, 1'b0, 0, 0) c1081105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081105));
	wire w1121105;
	repeater #(4, 1'b0, 0, 0) c1121105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121105));
	wire w1161105;
	repeater #(4, 1'b0, 0, 0) c1161105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161105));
	wire w1201105;
	repeater #(4, 1'b0, 0, 0) c1201105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201105));
	wire w1241105;
	repeater #(4, 1'b0, 0, 0) c1241105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241105));
	wire w1281105;
	repeater #(4, 1'b0, 0, 0) c1281105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281105));
	wire w1321105;
	repeater #(4, 1'b0, 0, 0) c1321105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321105));
	wire w1081106;
	repeater #(4, 1'b0, 0, 0) c1081106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081106));
	wire w1121106;
	repeater #(4, 1'b0, 0, 0) c1121106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121106));
	wire w1161106;
	repeater #(4, 1'b0, 0, 0) c1161106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161106));
	wire w1201106;
	repeater #(4, 1'b0, 0, 0) c1201106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201106));
	wire w1241106;
	repeater #(4, 1'b0, 0, 0) c1241106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241106));
	wire w1281106;
	repeater #(4, 1'b0, 0, 0) c1281106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281106));
	wire w1321106;
	repeater #(4, 1'b0, 0, 0) c1321106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321106));
	wire w1081107;
	repeater #(4, 1'b0, 0, 0) c1081107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081107));
	wire w1121107;
	repeater #(4, 1'b0, 0, 0) c1121107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121107));
	wire w1161107;
	repeater #(4, 1'b0, 0, 0) c1161107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161107));
	wire w1201107;
	repeater #(4, 1'b0, 0, 0) c1201107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201107));
	wire w1241107;
	repeater #(4, 1'b0, 0, 0) c1241107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241107));
	wire w1281107;
	repeater #(4, 1'b0, 0, 0) c1281107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281107));
	wire w1321107;
	repeater #(4, 1'b0, 0, 0) c1321107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321107));
	wire w1081108;
	repeater #(4, 1'b0, 0, 0) c1081108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081108));
	wire w1121108;
	repeater #(4, 1'b0, 0, 0) c1121108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121108));
	wire w1161108;
	repeater #(4, 1'b0, 0, 0) c1161108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161108));
	wire w1201108;
	repeater #(4, 1'b0, 0, 0) c1201108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201108));
	wire w1241108;
	repeater #(4, 1'b0, 0, 0) c1241108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241108));
	wire w1281108;
	repeater #(4, 1'b0, 0, 0) c1281108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281108));
	wire w1321108;
	repeater #(4, 1'b0, 0, 0) c1321108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321108));
	wire w1081109;
	repeater #(4, 1'b0, 0, 0) c1081109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081109));
	wire w1121109;
	repeater #(4, 1'b0, 0, 0) c1121109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121109));
	wire w1161109;
	repeater #(4, 1'b0, 0, 0) c1161109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161109));
	wire w1201109;
	repeater #(4, 1'b0, 0, 0) c1201109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201109));
	wire w1241109;
	repeater #(4, 1'b0, 0, 0) c1241109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241109));
	wire w1281109;
	repeater #(4, 1'b0, 0, 0) c1281109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281109));
	wire w1321109;
	repeater #(4, 1'b0, 0, 0) c1321109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321109));
	wire w1081110;
	repeater #(4, 1'b0, 0, 0) c1081110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081110));
	wire w1121110;
	repeater #(4, 1'b0, 0, 0) c1121110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121110));
	wire w1161110;
	repeater #(4, 1'b0, 0, 0) c1161110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161110));
	wire w1201110;
	repeater #(4, 1'b0, 0, 0) c1201110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201110));
	wire w1241110;
	repeater #(4, 1'b0, 0, 0) c1241110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241110));
	wire w1281110;
	repeater #(4, 1'b0, 0, 0) c1281110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281110));
	wire w1321110;
	repeater #(4, 1'b0, 0, 0) c1321110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321110));
	wire w1081111;
	repeater #(4, 1'b0, 0, 0) c1081111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081111));
	wire w1121111;
	repeater #(4, 1'b0, 0, 0) c1121111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121111));
	wire w1161111;
	repeater #(4, 1'b0, 0, 0) c1161111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161111));
	wire w1201111;
	repeater #(4, 1'b0, 0, 0) c1201111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201111));
	wire w1241111;
	repeater #(4, 1'b0, 0, 0) c1241111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241111));
	wire w1281111;
	repeater #(4, 1'b0, 0, 0) c1281111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281111));
	wire w1321111;
	repeater #(4, 1'b0, 0, 0) c1321111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321111));
	wire w1081112;
	repeater #(4, 1'b0, 0, 0) c1081112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081112));
	wire w1121112;
	repeater #(4, 1'b0, 0, 0) c1121112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121112));
	wire w1161112;
	repeater #(4, 1'b0, 0, 0) c1161112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161112));
	wire w1201112;
	repeater #(4, 1'b0, 0, 0) c1201112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201112));
	wire w1241112;
	repeater #(4, 1'b0, 0, 0) c1241112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241112));
	wire w1281112;
	repeater #(4, 1'b0, 0, 0) c1281112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281112));
	wire w1321112;
	repeater #(4, 1'b0, 0, 0) c1321112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321112));
	wire w1081113;
	repeater #(4, 1'b0, 0, 0) c1081113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081113));
	wire w1121113;
	repeater #(4, 1'b0, 0, 0) c1121113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121113));
	wire w1161113;
	repeater #(4, 1'b0, 0, 0) c1161113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161113));
	wire w1201113;
	repeater #(4, 1'b0, 0, 0) c1201113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201113));
	wire w1241113;
	repeater #(4, 1'b0, 0, 0) c1241113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241113));
	wire w1281113;
	repeater #(4, 1'b0, 0, 0) c1281113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281113));
	wire w1321113;
	repeater #(4, 1'b0, 0, 0) c1321113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321113));
	wire w1081114;
	repeater #(4, 1'b0, 0, 0) c1081114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081114));
	wire w1121114;
	repeater #(4, 1'b0, 0, 0) c1121114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121114));
	wire w1161114;
	repeater #(4, 1'b0, 0, 0) c1161114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161114));
	wire w1201114;
	repeater #(4, 1'b0, 0, 0) c1201114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201114));
	wire w1241114;
	repeater #(4, 1'b0, 0, 0) c1241114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241114));
	wire w1281114;
	repeater #(4, 1'b0, 0, 0) c1281114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281114));
	wire w1321114;
	repeater #(4, 1'b0, 0, 0) c1321114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321114));
	wire w1081115;
	repeater #(4, 1'b0, 0, 0) c1081115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081115));
	wire w1121115;
	repeater #(4, 1'b0, 0, 0) c1121115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121115));
	wire w1161115;
	repeater #(4, 1'b0, 0, 0) c1161115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161115));
	wire w1201115;
	repeater #(4, 1'b0, 0, 0) c1201115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201115));
	wire w1241115;
	repeater #(4, 1'b0, 0, 0) c1241115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241115));
	wire w1281115;
	repeater #(4, 1'b0, 0, 0) c1281115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281115));
	wire w1321115;
	repeater #(4, 1'b0, 0, 0) c1321115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321115));
	wire w1081116;
	repeater #(4, 1'b0, 0, 0) c1081116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081116));
	wire w1121116;
	repeater #(4, 1'b0, 0, 0) c1121116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121116));
	wire w1161116;
	repeater #(4, 1'b0, 0, 0) c1161116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161116));
	wire w1201116;
	repeater #(4, 1'b0, 0, 0) c1201116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201116));
	wire w1241116;
	repeater #(4, 1'b0, 0, 0) c1241116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241116));
	wire w1281116;
	repeater #(4, 1'b0, 0, 0) c1281116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281116));
	wire w1321116;
	repeater #(4, 1'b0, 0, 0) c1321116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321116));
	wire w1081117;
	repeater #(4, 1'b0, 0, 0) c1081117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081117));
	wire w1121117;
	repeater #(4, 1'b0, 0, 0) c1121117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121117));
	wire w1161117;
	repeater #(4, 1'b0, 0, 0) c1161117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161117));
	wire w1201117;
	repeater #(4, 1'b0, 0, 0) c1201117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201117));
	wire w1241117;
	repeater #(4, 1'b0, 0, 0) c1241117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241117));
	wire w1281117;
	repeater #(4, 1'b0, 0, 0) c1281117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281117));
	wire w1321117;
	repeater #(4, 1'b0, 0, 0) c1321117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321117));
	wire w1081118;
	repeater #(4, 1'b0, 0, 0) c1081118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081118));
	wire w1121118;
	repeater #(4, 1'b0, 0, 0) c1121118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121118));
	wire w1161118;
	repeater #(4, 1'b0, 0, 0) c1161118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161118));
	wire w1201118;
	repeater #(4, 1'b0, 0, 0) c1201118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201118));
	wire w1241118;
	repeater #(4, 1'b0, 0, 0) c1241118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241118));
	wire w1281118;
	repeater #(4, 1'b0, 0, 0) c1281118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281118));
	wire w1321118;
	repeater #(4, 1'b0, 0, 0) c1321118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321118));
	wire w1071126;
	repeater #(2, 1'b1, 0, 0) c1071126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1071126));
	wire w1081126;
	repeater #(1, 1'b0, 0, 0) c1081126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081126));
	wire w1111126;
	repeater #(2, 1'b1, 0, 0) c1111126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1111126));
	wire w1121126;
	repeater #(1, 1'b0, 0, 0) c1121126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121126));
	wire w1151126;
	repeater #(2, 1'b1, 0, 0) c1151126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1151126));
	wire w1161126;
	repeater #(1, 1'b0, 0, 0) c1161126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161126));
	wire w1191126;
	repeater #(2, 1'b1, 0, 0) c1191126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1191126));
	wire w1201126;
	repeater #(1, 1'b0, 0, 0) c1201126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201126));
	wire w1231126;
	repeater #(2, 1'b1, 0, 0) c1231126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1231126));
	wire w1241126;
	repeater #(1, 1'b0, 0, 0) c1241126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241126));
	wire w1271126;
	repeater #(2, 1'b1, 0, 0) c1271126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1271126));
	wire w1281126;
	repeater #(1, 1'b0, 0, 0) c1281126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281126));
	wire w1311126;
	repeater #(2, 1'b1, 0, 0) c1311126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1311126));
	wire w1321126;
	repeater #(1, 1'b0, 0, 0) c1321126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321126));
	wire w1071127;
	torch #(1'b0) c1071127 (.i_clk(tick), .i_in(), .o_out(w1071127));
	wire w1111127;
	torch #(1'b0) c1111127 (.i_clk(tick), .i_in(), .o_out(w1111127));
	wire w1151127;
	torch #(1'b0) c1151127 (.i_clk(tick), .i_in(), .o_out(w1151127));
	wire w1191127;
	torch #(1'b0) c1191127 (.i_clk(tick), .i_in(), .o_out(w1191127));
	wire w1231127;
	torch #(1'b0) c1231127 (.i_clk(tick), .i_in(), .o_out(w1231127));
	wire w1271127;
	torch #(1'b0) c1271127 (.i_clk(tick), .i_in(), .o_out(w1271127));
	wire w1311127;
	torch #(1'b0) c1311127 (.i_clk(tick), .i_in(), .o_out(w1311127));
	wire w1081128;
	repeater #(2, 1'b0, 0, 0) c1081128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081128));
	wire w1121128;
	repeater #(2, 1'b0, 0, 0) c1121128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121128));
	wire w1161128;
	repeater #(2, 1'b0, 0, 0) c1161128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161128));
	wire w1201128;
	repeater #(2, 1'b0, 0, 0) c1201128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201128));
	wire w1241128;
	repeater #(2, 1'b0, 0, 0) c1241128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241128));
	wire w1281128;
	repeater #(2, 1'b0, 0, 0) c1281128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281128));
	wire w1321128;
	repeater #(2, 1'b0, 0, 0) c1321128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321128));
	wire w1081129;
	repeater #(4, 1'b0, 0, 0) c1081129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081129));
	wire w1121129;
	repeater #(4, 1'b0, 0, 0) c1121129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121129));
	wire w1161129;
	repeater #(4, 1'b0, 0, 0) c1161129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161129));
	wire w1201129;
	repeater #(4, 1'b0, 0, 0) c1201129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201129));
	wire w1241129;
	repeater #(4, 1'b0, 0, 0) c1241129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241129));
	wire w1281129;
	repeater #(4, 1'b0, 0, 0) c1281129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281129));
	wire w1321129;
	repeater #(4, 1'b0, 0, 0) c1321129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321129));
	wire w1081130;
	repeater #(4, 1'b0, 0, 0) c1081130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081130));
	wire w1121130;
	repeater #(4, 1'b0, 0, 0) c1121130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121130));
	wire w1161130;
	repeater #(4, 1'b0, 0, 0) c1161130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161130));
	wire w1201130;
	repeater #(4, 1'b0, 0, 0) c1201130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201130));
	wire w1241130;
	repeater #(4, 1'b0, 0, 0) c1241130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241130));
	wire w1281130;
	repeater #(4, 1'b0, 0, 0) c1281130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281130));
	wire w1321130;
	repeater #(4, 1'b0, 0, 0) c1321130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321130));
	wire w1081131;
	repeater #(4, 1'b0, 0, 0) c1081131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081131));
	wire w1121131;
	repeater #(4, 1'b0, 0, 0) c1121131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121131));
	wire w1161131;
	repeater #(4, 1'b0, 0, 0) c1161131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161131));
	wire w1201131;
	repeater #(4, 1'b0, 0, 0) c1201131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201131));
	wire w1241131;
	repeater #(4, 1'b0, 0, 0) c1241131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241131));
	wire w1281131;
	repeater #(4, 1'b0, 0, 0) c1281131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281131));
	wire w1321131;
	repeater #(4, 1'b0, 0, 0) c1321131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321131));
	wire w1081132;
	repeater #(4, 1'b0, 0, 0) c1081132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081132));
	wire w1121132;
	repeater #(4, 1'b0, 0, 0) c1121132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121132));
	wire w1161132;
	repeater #(4, 1'b0, 0, 0) c1161132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161132));
	wire w1201132;
	repeater #(4, 1'b0, 0, 0) c1201132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201132));
	wire w1241132;
	repeater #(4, 1'b0, 0, 0) c1241132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241132));
	wire w1281132;
	repeater #(4, 1'b0, 0, 0) c1281132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281132));
	wire w1321132;
	repeater #(4, 1'b0, 0, 0) c1321132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321132));
	wire w1081133;
	repeater #(4, 1'b0, 0, 0) c1081133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081133));
	wire w1121133;
	repeater #(4, 1'b0, 0, 0) c1121133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121133));
	wire w1161133;
	repeater #(4, 1'b0, 0, 0) c1161133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161133));
	wire w1201133;
	repeater #(4, 1'b0, 0, 0) c1201133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201133));
	wire w1241133;
	repeater #(4, 1'b0, 0, 0) c1241133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241133));
	wire w1281133;
	repeater #(4, 1'b0, 0, 0) c1281133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281133));
	wire w1321133;
	repeater #(4, 1'b0, 0, 0) c1321133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321133));
	wire w1081134;
	repeater #(4, 1'b0, 0, 0) c1081134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081134));
	wire w1121134;
	repeater #(4, 1'b0, 0, 0) c1121134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121134));
	wire w1161134;
	repeater #(4, 1'b0, 0, 0) c1161134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161134));
	wire w1201134;
	repeater #(4, 1'b0, 0, 0) c1201134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201134));
	wire w1241134;
	repeater #(4, 1'b0, 0, 0) c1241134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241134));
	wire w1281134;
	repeater #(4, 1'b0, 0, 0) c1281134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281134));
	wire w1321134;
	repeater #(4, 1'b0, 0, 0) c1321134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321134));
	wire w1081135;
	repeater #(4, 1'b0, 0, 0) c1081135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081135));
	wire w1121135;
	repeater #(4, 1'b0, 0, 0) c1121135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1121135));
	wire w1161135;
	repeater #(4, 1'b0, 0, 0) c1161135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1161135));
	wire w1201135;
	repeater #(4, 1'b0, 0, 0) c1201135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201135));
	wire w1241135;
	repeater #(4, 1'b0, 0, 0) c1241135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1241135));
	wire w1281135;
	repeater #(4, 1'b0, 0, 0) c1281135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1281135));
	wire w1321135;
	repeater #(4, 1'b0, 0, 0) c1321135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1321135));
	wire w9200;
	repeater #(4, 1'b0, 0, 0) c9200 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9200));
	wire w9600;
	repeater #(4, 1'b0, 0, 0) c9600 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9600));
	wire w10000;
	repeater #(4, 1'b0, 0, 0) c10000 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10000));
	wire w10400;
	repeater #(4, 1'b0, 0, 0) c10400 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10400));
	wire w10800;
	repeater #(4, 1'b0, 0, 0) c10800 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10800));
	wire w11200;
	repeater #(4, 1'b0, 0, 0) c11200 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11200));
	wire w11600;
	repeater #(4, 1'b0, 0, 0) c11600 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11600));
	wire w9201;
	repeater #(4, 1'b0, 0, 0) c9201 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9201));
	wire w9601;
	repeater #(4, 1'b0, 0, 0) c9601 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9601));
	wire w10001;
	repeater #(4, 1'b0, 0, 0) c10001 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10001));
	wire w10401;
	repeater #(4, 1'b0, 0, 0) c10401 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10401));
	wire w10801;
	repeater #(4, 1'b0, 0, 0) c10801 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10801));
	wire w11201;
	repeater #(4, 1'b0, 0, 0) c11201 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11201));
	wire w11601;
	repeater #(4, 1'b0, 0, 0) c11601 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11601));
	wire w9202;
	repeater #(4, 1'b0, 0, 0) c9202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9202));
	wire w9602;
	repeater #(4, 1'b0, 0, 0) c9602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9602));
	wire w10002;
	repeater #(4, 1'b0, 0, 0) c10002 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10002));
	wire w10402;
	repeater #(4, 1'b0, 0, 0) c10402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10402));
	wire w10802;
	repeater #(4, 1'b0, 0, 0) c10802 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10802));
	wire w11202;
	repeater #(4, 1'b0, 0, 0) c11202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11202));
	wire w11602;
	repeater #(4, 1'b0, 0, 0) c11602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11602));
	wire w9203;
	repeater #(4, 1'b0, 0, 0) c9203 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9203));
	wire w9603;
	repeater #(4, 1'b0, 0, 0) c9603 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9603));
	wire w10003;
	repeater #(4, 1'b0, 0, 0) c10003 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10003));
	wire w10403;
	repeater #(4, 1'b0, 0, 0) c10403 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10403));
	wire w10803;
	repeater #(4, 1'b0, 0, 0) c10803 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10803));
	wire w11203;
	repeater #(4, 1'b0, 0, 0) c11203 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11203));
	wire w11603;
	repeater #(4, 1'b0, 0, 0) c11603 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11603));
	wire w9204;
	repeater #(4, 1'b0, 0, 0) c9204 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9204));
	wire w9604;
	repeater #(4, 1'b0, 0, 0) c9604 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9604));
	wire w10004;
	repeater #(4, 1'b0, 0, 0) c10004 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10004));
	wire w10404;
	repeater #(4, 1'b0, 0, 0) c10404 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10404));
	wire w10804;
	repeater #(4, 1'b0, 0, 0) c10804 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10804));
	wire w11204;
	repeater #(4, 1'b0, 0, 0) c11204 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11204));
	wire w11604;
	repeater #(4, 1'b0, 0, 0) c11604 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11604));
	wire w9205;
	repeater #(4, 1'b0, 0, 0) c9205 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9205));
	wire w9605;
	repeater #(4, 1'b0, 0, 0) c9605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9605));
	wire w10005;
	repeater #(4, 1'b0, 0, 0) c10005 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10005));
	wire w10405;
	repeater #(4, 1'b0, 0, 0) c10405 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10405));
	wire w10805;
	repeater #(4, 1'b0, 0, 0) c10805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10805));
	wire w11205;
	repeater #(4, 1'b0, 0, 0) c11205 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11205));
	wire w11605;
	repeater #(4, 1'b0, 0, 0) c11605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11605));
	wire w9206;
	repeater #(4, 1'b0, 0, 0) c9206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9206));
	wire w9606;
	repeater #(4, 1'b0, 0, 0) c9606 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9606));
	wire w10006;
	repeater #(4, 1'b0, 0, 0) c10006 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10006));
	wire w10406;
	repeater #(4, 1'b0, 0, 0) c10406 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10406));
	wire w10806;
	repeater #(4, 1'b0, 0, 0) c10806 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10806));
	wire w11206;
	repeater #(4, 1'b0, 0, 0) c11206 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11206));
	wire w11606;
	repeater #(4, 1'b0, 0, 0) c11606 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11606));
	wire w9207;
	repeater #(4, 1'b0, 0, 0) c9207 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9207));
	wire w9607;
	repeater #(4, 1'b0, 0, 0) c9607 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9607));
	wire w10007;
	repeater #(4, 1'b0, 0, 0) c10007 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10007));
	wire w10407;
	repeater #(4, 1'b0, 0, 0) c10407 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10407));
	wire w10807;
	repeater #(4, 1'b0, 0, 0) c10807 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10807));
	wire w11207;
	repeater #(4, 1'b0, 0, 0) c11207 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11207));
	wire w11607;
	repeater #(4, 1'b0, 0, 0) c11607 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11607));
	wire w121028;
	assign outputs[117] = ();
	wire w75065;
	torch #(1'b0) c75065 (.i_clk(tick), .i_in(), .o_out(w75065));
	wire w50092;
	repeater #(1, 1'b1, 0, 0) c50092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50092));
	wire w121124;
	repeater #(1, 1'b0, 0, 0) c121124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121124));
	wire w123124;

	wire w124124;
	repeater #(4, 1'b0, 0, 0) c124124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124124));
	wire w123125;
	repeater #(1, 1'b0, 0, 0) c123125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123125));
	wire w124126;
	repeater #(4, 1'b0, 0, 0) c124126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124126));
	wire w76165;
	repeater #(1, 1'b0, 0, 0) c76165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76165));
	wire w78165;
	repeater #(2, 1'b0, 0, 0) c78165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78165));
	wire w90168;
	repeater #(1, 1'b0, 0, 0) c90168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90168));
	wire w98168;
	repeater #(1, 1'b0, 0, 0) c98168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98168));
	wire w106168;
	repeater #(1, 1'b0, 0, 0) c106168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106168));
	wire w114168;
	repeater #(1, 1'b0, 0, 0) c114168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114168));
	wire w83169;
	repeater #(2, 1'b0, 0, 0) c83169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83169));
	wire w85169;
	repeater #(2, 1'b0, 0, 0) c85169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85169));
	wire w94169;
	repeater #(1, 1'b0, 0, 0) c94169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94169));
	wire w102169;
	repeater #(1, 1'b0, 0, 0) c102169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102169));
	wire w110169;
	repeater #(1, 1'b0, 0, 0) c110169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110169));
	wire w83170;
	repeater #(2, 1'b0, 0, 0) c83170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83170));
	wire w85170;
	repeater #(2, 1'b0, 0, 0) c85170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85170));
	wire w83171;
	repeater #(2, 1'b0, 0, 0) c83171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83171));
	wire w85171;
	repeater #(2, 1'b0, 0, 0) c85171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85171));
	wire w83172;
	repeater #(2, 1'b0, 0, 0) c83172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83172));
	wire w85172;
	repeater #(2, 1'b0, 0, 0) c85172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85172));
	wire w90172;
	torch #(1'b1) c90172 (.i_clk(tick), .i_in(), .o_out(w90172));
	wire w94172;
	torch #(1'b1) c94172 (.i_clk(tick), .i_in(), .o_out(w94172));
	wire w98172;
	torch #(1'b1) c98172 (.i_clk(tick), .i_in(), .o_out(w98172));
	wire w102172;
	torch #(1'b1) c102172 (.i_clk(tick), .i_in(), .o_out(w102172));
	wire w106172;
	torch #(1'b1) c106172 (.i_clk(tick), .i_in(), .o_out(w106172));
	wire w110172;
	torch #(1'b1) c110172 (.i_clk(tick), .i_in(), .o_out(w110172));
	wire w114172;
	torch #(1'b1) c114172 (.i_clk(tick), .i_in(), .o_out(w114172));
	wire w83173;
	repeater #(1, 1'b0, 0, 0) c83173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83173));
	wire w85173;
	repeater #(1, 1'b0, 0, 0) c85173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85173));
	wire w87175;
	repeater #(1, 1'b0, 0, 0) c87175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87175));
	wire w87176;
	repeater #(2, 1'b0, 0, 0) c87176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87176));
	wire w87177;
	repeater #(2, 1'b0, 0, 0) c87177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87177));
	wire w87178;
	repeater #(2, 1'b0, 0, 0) c87178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87178));
	wire w87179;
	repeater #(2, 1'b0, 0, 0) c87179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87179));
	wire w90187;
	torch #(1'b0) c90187 (.i_clk(tick), .i_in(), .o_out(w90187));
	wire w94187;
	torch #(1'b0) c94187 (.i_clk(tick), .i_in(), .o_out(w94187));
	wire w98187;
	torch #(1'b0) c98187 (.i_clk(tick), .i_in(), .o_out(w98187));
	wire w102187;
	torch #(1'b0) c102187 (.i_clk(tick), .i_in(), .o_out(w102187));
	wire w106187;
	torch #(1'b0) c106187 (.i_clk(tick), .i_in(), .o_out(w106187));
	wire w110187;
	torch #(1'b0) c110187 (.i_clk(tick), .i_in(), .o_out(w110187));
	wire w114187;
	torch #(1'b0) c114187 (.i_clk(tick), .i_in(), .o_out(w114187));
	wire w49191;

	wire w90192;
	repeater #(1, 1'b0, 0, 0) c90192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90192));
	wire w98192;
	repeater #(1, 1'b0, 0, 0) c98192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98192));
	wire w106192;
	repeater #(1, 1'b0, 0, 0) c106192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w106192));
	wire w114192;
	repeater #(1, 1'b0, 0, 0) c114192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w114192));
	wire w94193;
	repeater #(1, 1'b0, 0, 0) c94193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94193));
	wire w102193;
	repeater #(1, 1'b0, 0, 0) c102193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w102193));
	wire w110193;
	repeater #(1, 1'b0, 0, 0) c110193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110193));
	wire w90196;
	torch #(1'b1) c90196 (.i_clk(tick), .i_in(), .o_out(w90196));
	wire w94196;
	torch #(1'b1) c94196 (.i_clk(tick), .i_in(), .o_out(w94196));
	wire w98196;
	torch #(1'b1) c98196 (.i_clk(tick), .i_in(), .o_out(w98196));
	wire w102196;
	torch #(1'b1) c102196 (.i_clk(tick), .i_in(), .o_out(w102196));
	wire w106196;
	torch #(1'b1) c106196 (.i_clk(tick), .i_in(), .o_out(w106196));
	wire w110196;
	torch #(1'b1) c110196 (.i_clk(tick), .i_in(), .o_out(w110196));
	wire w114196;
	torch #(1'b1) c114196 (.i_clk(tick), .i_in(), .o_out(w114196));
	wire w901111;
	torch #(1'b0) c901111 (.i_clk(tick), .i_in(), .o_out(w901111));
	wire w941111;
	torch #(1'b0) c941111 (.i_clk(tick), .i_in(), .o_out(w941111));
	wire w981111;
	torch #(1'b0) c981111 (.i_clk(tick), .i_in(), .o_out(w981111));
	wire w1021111;
	torch #(1'b0) c1021111 (.i_clk(tick), .i_in(), .o_out(w1021111));
	wire w1061111;
	torch #(1'b0) c1061111 (.i_clk(tick), .i_in(), .o_out(w1061111));
	wire w1101111;
	torch #(1'b0) c1101111 (.i_clk(tick), .i_in(), .o_out(w1101111));
	wire w1141111;
	torch #(1'b0) c1141111 (.i_clk(tick), .i_in(), .o_out(w1141111));
	wire w1911114;
	repeater #(1, 1'b0, 0, 0) c1911114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911114));
	wire w901116;
	repeater #(1, 1'b0, 0, 0) c901116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901116));
	wire w981116;
	repeater #(1, 1'b0, 0, 0) c981116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981116));
	wire w1061116;
	repeater #(1, 1'b0, 0, 0) c1061116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061116));
	wire w1141116;
	repeater #(1, 1'b0, 0, 0) c1141116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1141116));
	wire w941117;
	repeater #(1, 1'b0, 0, 0) c941117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941117));
	wire w1021117;
	repeater #(1, 1'b0, 0, 0) c1021117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1021117));
	wire w1101117;
	repeater #(1, 1'b0, 0, 0) c1101117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101117));
	wire w901120;
	torch #(1'b1) c901120 (.i_clk(tick), .i_in(), .o_out(w901120));
	wire w941120;
	torch #(1'b1) c941120 (.i_clk(tick), .i_in(), .o_out(w941120));
	wire w981120;
	torch #(1'b1) c981120 (.i_clk(tick), .i_in(), .o_out(w981120));
	wire w1021120;
	torch #(1'b1) c1021120 (.i_clk(tick), .i_in(), .o_out(w1021120));
	wire w1061120;
	torch #(1'b1) c1061120 (.i_clk(tick), .i_in(), .o_out(w1061120));
	wire w1101120;
	torch #(1'b1) c1101120 (.i_clk(tick), .i_in(), .o_out(w1101120));
	wire w1141120;
	torch #(1'b1) c1141120 (.i_clk(tick), .i_in(), .o_out(w1141120));
	wire w901135;
	torch #(1'b0) c901135 (.i_clk(tick), .i_in(), .o_out(w901135));
	wire w941135;
	torch #(1'b0) c941135 (.i_clk(tick), .i_in(), .o_out(w941135));
	wire w981135;
	torch #(1'b0) c981135 (.i_clk(tick), .i_in(), .o_out(w981135));
	wire w1021135;
	torch #(1'b0) c1021135 (.i_clk(tick), .i_in(), .o_out(w1021135));
	wire w1061135;
	torch #(1'b0) c1061135 (.i_clk(tick), .i_in(), .o_out(w1061135));
	wire w1101135;
	torch #(1'b0) c1101135 (.i_clk(tick), .i_in(), .o_out(w1101135));
	wire w1141135;
	torch #(1'b0) c1141135 (.i_clk(tick), .i_in(), .o_out(w1141135));
	wire w7404;
	repeater #(1, 1'b0, 0, 0) c7404 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7404));
	wire w8204;
	repeater #(1, 1'b0, 0, 0) c8204 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8204));
	wire w9004;
	repeater #(1, 1'b0, 0, 0) c9004 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9004));
	wire w9804;
	repeater #(1, 1'b0, 0, 0) c9804 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9804));
	wire w7805;
	repeater #(1, 1'b0, 0, 0) c7805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7805));
	wire w8605;
	repeater #(1, 1'b0, 0, 0) c8605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8605));
	wire w9405;
	repeater #(1, 1'b0, 0, 0) c9405 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9405));
	wire w7408;
	torch #(1'b1) c7408 (.i_clk(tick), .i_in(), .o_out(w7408));
	wire w7808;
	torch #(1'b1) c7808 (.i_clk(tick), .i_in(), .o_out(w7808));
	wire w8208;
	torch #(1'b1) c8208 (.i_clk(tick), .i_in(), .o_out(w8208));
	wire w8608;
	torch #(1'b1) c8608 (.i_clk(tick), .i_in(), .o_out(w8608));
	wire w9008;
	torch #(1'b1) c9008 (.i_clk(tick), .i_in(), .o_out(w9008));
	wire w9408;
	torch #(1'b1) c9408 (.i_clk(tick), .i_in(), .o_out(w9408));
	wire w9808;
	torch #(1'b1) c9808 (.i_clk(tick), .i_in(), .o_out(w9808));
	wire w74023;
	torch #(1'b0) c74023 (.i_clk(tick), .i_in(), .o_out(w74023));
	wire w78023;
	torch #(1'b0) c78023 (.i_clk(tick), .i_in(), .o_out(w78023));
	wire w82023;
	torch #(1'b0) c82023 (.i_clk(tick), .i_in(), .o_out(w82023));
	wire w86023;
	torch #(1'b0) c86023 (.i_clk(tick), .i_in(), .o_out(w86023));
	wire w90023;
	torch #(1'b0) c90023 (.i_clk(tick), .i_in(), .o_out(w90023));
	wire w94023;
	torch #(1'b0) c94023 (.i_clk(tick), .i_in(), .o_out(w94023));
	wire w98023;
	torch #(1'b0) c98023 (.i_clk(tick), .i_in(), .o_out(w98023));
	wire w74028;
	repeater #(1, 1'b0, 0, 0) c74028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74028));
	wire w82028;
	repeater #(1, 1'b0, 0, 0) c82028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82028));
	wire w90028;
	repeater #(1, 1'b0, 0, 0) c90028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90028));
	wire w98028;
	repeater #(1, 1'b0, 0, 0) c98028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98028));
	wire w78029;
	repeater #(1, 1'b0, 0, 0) c78029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78029));
	wire w86029;
	repeater #(1, 1'b0, 0, 0) c86029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86029));
	wire w94029;
	repeater #(1, 1'b0, 0, 0) c94029 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94029));
	wire w74032;
	torch #(1'b1) c74032 (.i_clk(tick), .i_in(), .o_out(w74032));
	wire w78032;
	torch #(1'b1) c78032 (.i_clk(tick), .i_in(), .o_out(w78032));
	wire w82032;
	torch #(1'b1) c82032 (.i_clk(tick), .i_in(), .o_out(w82032));
	wire w86032;
	torch #(1'b1) c86032 (.i_clk(tick), .i_in(), .o_out(w86032));
	wire w90032;
	torch #(1'b1) c90032 (.i_clk(tick), .i_in(), .o_out(w90032));
	wire w94032;
	torch #(1'b1) c94032 (.i_clk(tick), .i_in(), .o_out(w94032));
	wire w98032;
	torch #(1'b1) c98032 (.i_clk(tick), .i_in(), .o_out(w98032));
	wire w74047;
	torch #(1'b0) c74047 (.i_clk(tick), .i_in(), .o_out(w74047));
	wire w78047;
	torch #(1'b0) c78047 (.i_clk(tick), .i_in(), .o_out(w78047));
	wire w82047;
	torch #(1'b0) c82047 (.i_clk(tick), .i_in(), .o_out(w82047));
	wire w86047;
	torch #(1'b0) c86047 (.i_clk(tick), .i_in(), .o_out(w86047));
	wire w90047;
	torch #(1'b0) c90047 (.i_clk(tick), .i_in(), .o_out(w90047));
	wire w94047;
	torch #(1'b0) c94047 (.i_clk(tick), .i_in(), .o_out(w94047));
	wire w98047;
	torch #(1'b0) c98047 (.i_clk(tick), .i_in(), .o_out(w98047));
	wire w600104;
	repeater #(1, 1'b0, 0, 0) c600104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w600104));
	wire w530106;
	repeater #(1, 1'b0, 0, 0) c530106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w530106));
	wire w550106;

	wire w670106;
	repeater #(2, 1'b0, 0, 0) c670106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w670106));
	wire w660107;
	repeater #(2, 1'b0, 0, 0) c660107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660107));
	wire w680107;
	repeater #(2, 1'b0, 0, 0) c680107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w680107));
	wire w1790107;
	repeater #(1, 1'b0, 0, 0) c1790107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1790107));
	wire w1970107;
	repeater #(1, 1'b0, 0, 0) c1970107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1970107));
	wire w70108;
	repeater #(1, 1'b0, 0, 0) c70108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70108));
	wire w250108;
	repeater #(1, 1'b0, 0, 0) c250108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w250108));
	wire w430108;
	repeater #(1, 1'b0, 0, 0) c430108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w430108));
	wire w580108;

	wire w640108;
	repeater #(1, 1'b0, 0, 0) c640108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w640108));
	wire w650108;
	repeater #(2, 1'b0, 0, 0) c650108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w650108));
	wire w1000108;
	torch #(1'b0) c1000108 (.i_clk(tick), .i_in(), .o_out(w1000108));
	wire w1030108;
	torch #(1'b1) c1030108 (.i_clk(tick), .i_in(), .o_out(w1030108));
	wire w1830109;
	repeater #(1, 1'b0, 0, 0) c1830109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1830109));
	wire w2010109;
	repeater #(1, 1'b0, 0, 0) c2010109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2010109));
	wire w110110;
	repeater #(1, 1'b0, 0, 0) c110110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110110));
	wire w290110;
	repeater #(1, 1'b0, 0, 0) c290110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w290110));
	wire w470110;
	repeater #(1, 1'b0, 0, 0) c470110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470110));
	wire w760113;
	repeater #(1, 1'b1, 0, 0) c760113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w760113));
	wire w800113;
	repeater #(1, 1'b1, 0, 0) c800113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800113));
	wire w840113;
	repeater #(1, 1'b1, 0, 0) c840113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840113));
	wire w880113;
	repeater #(1, 1'b1, 0, 0) c880113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w880113));
	wire w920113;
	repeater #(1, 1'b1, 0, 0) c920113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w920113));
	wire w960113;
	repeater #(1, 1'b1, 0, 0) c960113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w960113));
	wire w1000113;
	repeater #(1, 1'b1, 0, 0) c1000113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1000113));
	wire w340120;
	repeater #(1, 1'b1, 0, 0) c340120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340120));
	wire w1750121;
	repeater #(1, 1'b0, 0, 0) c1750121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750121));
	wire w1770121;
	repeater #(1, 1'b0, 0, 0) c1770121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770121));
	wire w1000132;
	torch #(1'b0) c1000132 (.i_clk(tick), .i_in(), .o_out(w1000132));
	wire w1030132;
	torch #(1'b1) c1030132 (.i_clk(tick), .i_in(), .o_out(w1030132));
	wire w1060133;
	repeater #(1, 1'b1, 0, 0) c1060133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060133));
	wire w1080133;
	repeater #(1, 1'b1, 0, 0) c1080133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1080133));
	wire w760137;
	repeater #(1, 1'b1, 0, 0) c760137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w760137));
	wire w800137;
	repeater #(1, 1'b1, 0, 0) c800137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800137));
	wire w840137;
	repeater #(1, 1'b1, 0, 0) c840137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840137));
	wire w880137;
	repeater #(1, 1'b1, 0, 0) c880137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w880137));
	wire w920137;
	repeater #(1, 1'b1, 0, 0) c920137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w920137));
	wire w960137;
	repeater #(1, 1'b1, 0, 0) c960137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w960137));
	wire w1000137;
	repeater #(1, 1'b1, 0, 0) c1000137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1000137));
	wire w1750139;
	repeater #(1, 1'b0, 0, 0) c1750139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1750139));
	wire w1770139;
	repeater #(1, 1'b0, 0, 0) c1770139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770139));
	wire w1060155;
	repeater #(1, 1'b1, 0, 0) c1060155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1060155));
	wire w1100155;
	repeater #(1, 1'b1, 0, 0) c1100155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1100155));
	wire w1000156;
	torch #(1'b0) c1000156 (.i_clk(tick), .i_in(), .o_out(w1000156));
	wire w1030156;
	torch #(1'b1) c1030156 (.i_clk(tick), .i_in(), .o_out(w1030156));
	wire w1770157;
	repeater #(1, 1'b0, 0, 0) c1770157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1770157));
	wire w760161;
	repeater #(1, 1'b1, 0, 0) c760161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w760161));
	wire w800161;
	repeater #(1, 1'b1, 0, 0) c800161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w800161));
	wire w840161;
	repeater #(1, 1'b1, 0, 0) c840161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840161));
	wire w880161;
	repeater #(1, 1'b1, 0, 0) c880161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w880161));
	wire w920161;
	repeater #(1, 1'b1, 0, 0) c920161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w920161));
	wire w960161;
	repeater #(1, 1'b1, 0, 0) c960161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w960161));
	wire w1000161;
	repeater #(1, 1'b1, 0, 0) c1000161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1000161));
	wire w10610;
	repeater #(1, 1'b1, 0, 0) c10610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10610));
	wire w10011;
	torch #(1'b0) c10011 (.i_clk(tick), .i_in(), .o_out(w10011));
	wire w10311;
	torch #(1'b1) c10311 (.i_clk(tick), .i_in(), .o_out(w10311));
	wire w7616;
	repeater #(1, 1'b1, 0, 0) c7616 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7616));
	wire w8016;
	repeater #(1, 1'b1, 0, 0) c8016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8016));
	wire w8416;
	repeater #(1, 1'b1, 0, 0) c8416 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8416));
	wire w8816;
	repeater #(1, 1'b1, 0, 0) c8816 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8816));
	wire w9216;
	repeater #(1, 1'b1, 0, 0) c9216 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9216));
	wire w9616;
	repeater #(1, 1'b1, 0, 0) c9616 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9616));
	wire w10016;
	repeater #(1, 1'b1, 0, 0) c10016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10016));
	wire w108124;
	repeater #(1, 1'b1, 0, 0) c108124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w108124));
	wire w110124;
	repeater #(1, 1'b1, 0, 0) c110124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w110124));
	wire w100125;
	torch #(1'b0) c100125 (.i_clk(tick), .i_in(), .o_out(w100125));
	wire w103125;
	torch #(1'b1) c103125 (.i_clk(tick), .i_in(), .o_out(w103125));
	wire w76130;
	repeater #(1, 1'b1, 0, 0) c76130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w76130));
	wire w80130;
	repeater #(1, 1'b1, 0, 0) c80130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80130));
	wire w84130;
	repeater #(1, 1'b1, 0, 0) c84130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84130));
	wire w88130;
	repeater #(1, 1'b1, 0, 0) c88130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88130));
	wire w92130;
	repeater #(1, 1'b1, 0, 0) c92130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92130));
	wire w96130;
	repeater #(1, 1'b1, 0, 0) c96130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w96130));
	wire w100130;
	repeater #(1, 1'b1, 0, 0) c100130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100130));
	wire w104148;
	torch #(1'b1) c104148 (.i_clk(tick), .i_in(), .o_out(w104148));
	wire w891107;
	repeater #(1, 1'b1, 0, 0) c891107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w891107));
	wire w1061109;
	repeater #(1, 1'b1, 0, 0) c1061109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061109));
	wire w1081109;
	repeater #(1, 1'b1, 0, 0) c1081109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1081109));
	wire w1101109;
	repeater #(1, 1'b1, 0, 0) c1101109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101109));
	wire w671111;
	repeater #(1, 1'b0, 0, 0) c671111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w671111));
	wire w691111;
	repeater #(1, 1'b0, 0, 0) c691111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691111));
	wire w741111;
	repeater #(1, 1'b0, 0, 0) c741111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741111));
	wire w751111;

	wire w781111;
	repeater #(1, 1'b0, 0, 0) c781111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w781111));
	wire w791111;

	wire w821111;
	repeater #(1, 1'b0, 0, 0) c821111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821111));
	wire w831111;

	wire w861111;
	repeater #(1, 1'b0, 0, 0) c861111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861111));
	wire w871111;

	wire w901111;
	repeater #(1, 1'b0, 0, 0) c901111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901111));
	wire w911111;

	wire w941111;
	repeater #(1, 1'b0, 0, 0) c941111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941111));
	wire w951111;

	wire w981111;
	repeater #(1, 1'b0, 0, 0) c981111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981111));
	wire w991111;

	wire w671112;
	repeater #(2, 1'b0, 0, 0) c671112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w671112));
	wire w691112;
	repeater #(2, 1'b0, 0, 0) c691112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691112));
	wire w671113;
	repeater #(2, 1'b0, 0, 0) c671113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w671113));
	wire w691113;
	repeater #(2, 1'b0, 0, 0) c691113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691113));
	wire w671114;
	repeater #(2, 1'b0, 0, 0) c671114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w671114));
	wire w691114;
	repeater #(2, 1'b0, 0, 0) c691114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691114));
	wire w741114;
	repeater #(1, 1'b0, 0, 0) c741114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741114));
	wire w791114;
	repeater #(1, 1'b0, 0, 0) c791114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791114));
	wire w821114;
	repeater #(1, 1'b0, 0, 0) c821114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821114));
	wire w871114;
	repeater #(1, 1'b0, 0, 0) c871114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w871114));
	wire w901114;
	repeater #(1, 1'b0, 0, 0) c901114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901114));
	wire w951114;
	repeater #(1, 1'b0, 0, 0) c951114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951114));
	wire w671115;
	repeater #(2, 1'b0, 0, 0) c671115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w671115));
	wire w691115;
	repeater #(2, 1'b0, 0, 0) c691115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w691115));
	wire w981115;
	repeater #(4, 1'b0, 0, 0) c981115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981115));
	wire w741116;
	repeater #(4, 1'b0, 0, 0) c741116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741116));
	wire w791116;
	repeater #(2, 1'b0, 0, 0) c791116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791116));
	wire w821116;
	repeater #(4, 1'b0, 0, 0) c821116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821116));
	wire w871116;
	repeater #(2, 1'b0, 0, 0) c871116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w871116));
	wire w901116;
	repeater #(4, 1'b0, 0, 0) c901116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901116));
	wire w951116;
	repeater #(2, 1'b0, 0, 0) c951116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951116));
	wire w791118;
	repeater #(2, 1'b0, 0, 0) c791118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791118));
	wire w871118;
	repeater #(2, 1'b0, 0, 0) c871118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w871118));
	wire w951118;
	repeater #(2, 1'b0, 0, 0) c951118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951118));
	wire w331119;

	wire w711119;
	repeater #(2, 1'b0, 0, 0) c711119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711119));
	wire w981119;
	repeater #(2, 1'b0, 0, 0) c981119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981119));
	wire w711120;
	repeater #(2, 1'b0, 0, 0) c711120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711120));
	wire w771120;
	repeater #(1, 1'b0, 0, 0) c771120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w771120));
	wire w851120;
	repeater #(1, 1'b1, 0, 0) c851120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w851120));
	wire w931120;
	repeater #(1, 1'b1, 0, 0) c931120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w931120));
	wire w711121;
	repeater #(2, 1'b0, 0, 0) c711121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711121));
	wire w741121;

	wire w751121;

	wire w791121;

	wire w821121;

	wire w831121;

	wire w871121;

	wire w901121;

	wire w911121;

	wire w951121;

	wire w711122;
	repeater #(2, 1'b0, 0, 0) c711122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711122));
	wire w711123;
	repeater #(1, 1'b0, 0, 0) c711123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w711123));
	wire w741124;
	repeater #(1, 1'b0, 0, 0) c741124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741124));
	wire w791124;
	repeater #(1, 1'b0, 0, 0) c791124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791124));
	wire w901124;
	repeater #(1, 1'b0, 0, 0) c901124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901124));
	wire w951124;
	repeater #(1, 1'b0, 0, 0) c951124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951124));
	wire w741126;
	repeater #(4, 1'b0, 0, 0) c741126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741126));
	wire w791126;
	repeater #(2, 1'b0, 0, 0) c791126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791126));
	wire w801126;
	repeater #(1, 1'b0, 0, 0) c801126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w801126));
	wire w821126;
	repeater #(4, 1'b0, 0, 0) c821126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821126));
	wire w901126;
	repeater #(4, 1'b0, 0, 0) c901126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901126));
	wire w951126;
	repeater #(2, 1'b0, 0, 0) c951126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951126));
	wire w821127;
	repeater #(1, 1'b0, 0, 0) c821127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821127));
	wire w861127;
	repeater #(3, 1'b0, 0, 0) c861127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861127));
	wire w791128;
	repeater #(2, 1'b0, 0, 0) c791128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w791128));
	wire w951128;
	repeater #(2, 1'b0, 0, 0) c951128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w951128));
	wire w871129;
	repeater #(1, 1'b0, 0, 0) c871129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w871129));
	wire w881129;
	repeater #(1, 1'b0, 0, 0) c881129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w881129));
	wire w771130;
	repeater #(1, 1'b0, 0, 0) c771130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w771130));
	wire w851130;
	repeater #(1, 1'b1, 0, 0) c851130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w851130));
	wire w871130;
	repeater #(4, 1'b0, 0, 0) c871130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w871130));
	wire w931130;
	repeater #(1, 1'b1, 0, 0) c931130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w931130));
	wire w741131;

	wire w751131;

	wire w791131;

	wire w821131;

	wire w831131;

	wire w871131;

	wire w901131;

	wire w911131;

	wire w951131;

	wire w1091132;
	torch #(1'b1) c1091132 (.i_clk(tick), .i_in(), .o_out(w1091132));
	wire w741135;
	repeater #(1, 1'b0, 0, 0) c741135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w741135));
	wire w751135;

	wire w781135;
	repeater #(1, 1'b0, 0, 0) c781135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w781135));
	wire w791135;

	wire w821135;
	repeater #(1, 1'b0, 0, 0) c821135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w821135));
	wire w831135;

	wire w861135;
	repeater #(1, 1'b0, 0, 0) c861135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w861135));
	wire w871135;

	wire w901135;
	repeater #(1, 1'b0, 0, 0) c901135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901135));
	wire w911135;

	wire w941135;
	repeater #(1, 1'b0, 0, 0) c941135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941135));
	wire w951135;

	wire w981135;
	repeater #(1, 1'b0, 0, 0) c981135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981135));
	wire w991135;

	wire w5802;
	repeater #(1, 1'b0, 0, 0) c5802 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5802));
	wire w6302;
	repeater #(1, 1'b0, 0, 0) c6302 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6302));
	wire w6602;
	repeater #(1, 1'b0, 0, 0) c6602 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6602));
	wire w7102;
	repeater #(1, 1'b0, 0, 0) c7102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7102));
	wire w7402;
	repeater #(1, 1'b0, 0, 0) c7402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7402));
	wire w7902;
	repeater #(1, 1'b0, 0, 0) c7902 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7902));
	wire w8203;
	repeater #(4, 1'b0, 0, 0) c8203 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8203));
	wire w5804;
	repeater #(4, 1'b0, 0, 0) c5804 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5804));
	wire w6304;
	repeater #(2, 1'b0, 0, 0) c6304 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6304));
	wire w6604;
	repeater #(4, 1'b0, 0, 0) c6604 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6604));
	wire w7104;
	repeater #(2, 1'b0, 0, 0) c7104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7104));
	wire w7404;
	repeater #(4, 1'b0, 0, 0) c7404 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7404));
	wire w7904;
	repeater #(2, 1'b0, 0, 0) c7904 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7904));
	wire w6306;
	repeater #(2, 1'b0, 0, 0) c6306 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6306));
	wire w7106;
	repeater #(2, 1'b0, 0, 0) c7106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7106));
	wire w7906;
	repeater #(2, 1'b0, 0, 0) c7906 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7906));
	wire w8207;
	repeater #(2, 1'b0, 0, 0) c8207 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8207));
	wire w6108;
	repeater #(1, 1'b1, 0, 0) c6108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6108));
	wire w6908;
	repeater #(1, 1'b0, 0, 0) c6908 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6908));
	wire w7708;
	repeater #(1, 1'b1, 0, 0) c7708 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7708));
	wire w5809;

	wire w5909;

	wire w6309;

	wire w6609;

	wire w6709;

	wire w7109;

	wire w7409;

	wire w7509;

	wire w7909;

	wire w58012;
	repeater #(1, 1'b0, 0, 0) c58012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58012));
	wire w63012;
	repeater #(1, 1'b0, 0, 0) c63012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63012));
	wire w74012;
	repeater #(1, 1'b0, 0, 0) c74012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74012));
	wire w79012;
	repeater #(1, 1'b0, 0, 0) c79012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79012));
	wire w58014;
	repeater #(4, 1'b0, 0, 0) c58014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58014));
	wire w63014;
	repeater #(2, 1'b0, 0, 0) c63014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63014));
	wire w64014;
	repeater #(1, 1'b0, 0, 0) c64014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64014));
	wire w66014;
	repeater #(4, 1'b0, 0, 0) c66014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66014));
	wire w74014;
	repeater #(4, 1'b0, 0, 0) c74014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74014));
	wire w79014;
	repeater #(2, 1'b0, 0, 0) c79014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79014));
	wire w66015;
	repeater #(1, 1'b0, 0, 0) c66015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66015));
	wire w70015;
	repeater #(3, 1'b0, 0, 0) c70015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70015));
	wire w63016;
	repeater #(2, 1'b0, 0, 0) c63016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63016));
	wire w79016;
	repeater #(2, 1'b0, 0, 0) c79016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79016));
	wire w71017;
	repeater #(1, 1'b0, 0, 0) c71017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71017));
	wire w72017;
	repeater #(1, 1'b0, 0, 0) c72017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72017));
	wire w61018;
	repeater #(1, 1'b0, 0, 0) c61018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61018));
	wire w69018;
	repeater #(1, 1'b1, 0, 0) c69018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69018));
	wire w71018;
	repeater #(4, 1'b0, 0, 0) c71018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71018));
	wire w77018;
	repeater #(1, 1'b1, 0, 0) c77018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77018));
	wire w58019;

	wire w59019;

	wire w63019;

	wire w66019;

	wire w67019;

	wire w71019;

	wire w74019;

	wire w75019;

	wire w79019;

	wire w91020;
	torch #(1'b1) c91020 (.i_clk(tick), .i_in(), .o_out(w91020));
	wire w58023;
	repeater #(1, 1'b0, 0, 0) c58023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58023));
	wire w59023;

	wire w62023;
	repeater #(1, 1'b0, 0, 0) c62023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62023));
	wire w63023;

	wire w66023;
	repeater #(1, 1'b0, 0, 0) c66023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66023));
	wire w67023;

	wire w70023;
	repeater #(1, 1'b0, 0, 0) c70023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70023));
	wire w71023;

	wire w74023;
	repeater #(1, 1'b0, 0, 0) c74023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74023));
	wire w75023;

	wire w78023;
	repeater #(1, 1'b0, 0, 0) c78023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78023));
	wire w79023;

	wire w82023;
	repeater #(1, 1'b0, 0, 0) c82023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82023));
	wire w83023;

	wire w58026;
	repeater #(1, 1'b0, 0, 0) c58026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58026));
	wire w63026;
	repeater #(1, 1'b0, 0, 0) c63026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63026));
	wire w66026;
	repeater #(1, 1'b0, 0, 0) c66026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66026));
	wire w71026;
	repeater #(1, 1'b0, 0, 0) c71026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71026));
	wire w74026;
	repeater #(1, 1'b0, 0, 0) c74026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74026));
	wire w79026;
	repeater #(1, 1'b0, 0, 0) c79026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79026));
	wire w82027;
	repeater #(4, 1'b0, 0, 0) c82027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82027));
	wire w58028;
	repeater #(4, 1'b0, 0, 0) c58028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58028));
	wire w63028;
	repeater #(2, 1'b0, 0, 0) c63028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63028));
	wire w66028;
	repeater #(4, 1'b0, 0, 0) c66028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66028));
	wire w71028;
	repeater #(2, 1'b0, 0, 0) c71028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71028));
	wire w74028;
	repeater #(4, 1'b0, 0, 0) c74028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74028));
	wire w79028;
	repeater #(2, 1'b0, 0, 0) c79028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79028));
	wire w63030;
	repeater #(2, 1'b0, 0, 0) c63030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63030));
	wire w71030;
	repeater #(2, 1'b0, 0, 0) c71030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71030));
	wire w79030;
	repeater #(2, 1'b0, 0, 0) c79030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79030));
	wire w82031;
	repeater #(2, 1'b0, 0, 0) c82031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82031));
	wire w61032;
	repeater #(1, 1'b0, 0, 0) c61032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61032));
	wire w69032;
	repeater #(1, 1'b0, 0, 0) c69032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69032));
	wire w77032;
	repeater #(1, 1'b1, 0, 0) c77032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77032));
	wire w58033;

	wire w59033;

	wire w63033;

	wire w66033;

	wire w67033;

	wire w71033;

	wire w74033;

	wire w75033;

	wire w79033;

	wire w58036;
	repeater #(1, 1'b0, 0, 0) c58036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58036));
	wire w63036;
	repeater #(1, 1'b0, 0, 0) c63036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63036));
	wire w74036;
	repeater #(1, 1'b0, 0, 0) c74036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74036));
	wire w79036;
	repeater #(1, 1'b0, 0, 0) c79036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79036));
	wire w58038;
	repeater #(4, 1'b0, 0, 0) c58038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58038));
	wire w63038;
	repeater #(2, 1'b0, 0, 0) c63038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63038));
	wire w64038;
	repeater #(1, 1'b0, 0, 0) c64038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64038));
	wire w66038;
	repeater #(4, 1'b0, 0, 0) c66038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66038));
	wire w74038;
	repeater #(4, 1'b0, 0, 0) c74038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74038));
	wire w79038;
	repeater #(2, 1'b0, 0, 0) c79038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79038));
	wire w66039;
	repeater #(1, 1'b0, 0, 0) c66039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66039));
	wire w70039;
	repeater #(3, 1'b0, 0, 0) c70039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70039));
	wire w63040;
	repeater #(2, 1'b0, 0, 0) c63040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63040));
	wire w79040;
	repeater #(2, 1'b0, 0, 0) c79040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79040));
	wire w71041;
	repeater #(1, 1'b0, 0, 0) c71041 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71041));
	wire w72041;
	repeater #(1, 1'b0, 0, 0) c72041 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72041));
	wire w61042;
	repeater #(1, 1'b0, 0, 0) c61042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61042));
	wire w69042;
	repeater #(1, 1'b1, 0, 0) c69042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69042));
	wire w71042;
	repeater #(4, 1'b0, 0, 0) c71042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71042));
	wire w77042;
	repeater #(1, 1'b1, 0, 0) c77042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77042));
	wire w58043;

	wire w59043;

	wire w63043;

	wire w66043;

	wire w67043;

	wire w71043;

	wire w74043;

	wire w75043;

	wire w79043;

	wire w91044;
	torch #(1'b1) c91044 (.i_clk(tick), .i_in(), .o_out(w91044));
	wire w93044;
	torch #(1'b1) c93044 (.i_clk(tick), .i_in(), .o_out(w93044));
	wire w58047;
	repeater #(1, 1'b0, 0, 0) c58047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58047));
	wire w59047;

	wire w62047;
	repeater #(1, 1'b0, 0, 0) c62047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62047));
	wire w63047;

	wire w66047;
	repeater #(1, 1'b0, 0, 0) c66047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66047));
	wire w67047;

	wire w70047;
	repeater #(1, 1'b0, 0, 0) c70047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70047));
	wire w71047;

	wire w74047;
	repeater #(1, 1'b0, 0, 0) c74047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74047));
	wire w75047;

	wire w78047;
	repeater #(1, 1'b0, 0, 0) c78047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78047));
	wire w79047;

	wire w82047;
	repeater #(1, 1'b0, 0, 0) c82047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82047));
	wire w83047;

	wire w58050;
	repeater #(1, 1'b0, 0, 0) c58050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58050));
	wire w63050;
	repeater #(1, 1'b0, 0, 0) c63050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63050));
	wire w66050;
	repeater #(1, 1'b0, 0, 0) c66050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66050));
	wire w71050;
	repeater #(1, 1'b0, 0, 0) c71050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71050));
	wire w74050;
	repeater #(1, 1'b0, 0, 0) c74050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74050));
	wire w79050;
	repeater #(1, 1'b0, 0, 0) c79050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79050));
	wire w82051;
	repeater #(4, 1'b0, 0, 0) c82051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82051));
	wire w58052;
	repeater #(4, 1'b0, 0, 0) c58052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58052));
	wire w63052;
	repeater #(2, 1'b0, 0, 0) c63052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63052));
	wire w66052;
	repeater #(4, 1'b0, 0, 0) c66052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66052));
	wire w71052;
	repeater #(2, 1'b0, 0, 0) c71052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71052));
	wire w74052;
	repeater #(4, 1'b0, 0, 0) c74052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74052));
	wire w79052;
	repeater #(2, 1'b0, 0, 0) c79052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79052));
	wire w63054;
	repeater #(2, 1'b0, 0, 0) c63054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63054));
	wire w71054;
	repeater #(2, 1'b0, 0, 0) c71054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71054));
	wire w79054;
	repeater #(2, 1'b0, 0, 0) c79054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79054));
	wire w82055;
	repeater #(2, 1'b0, 0, 0) c82055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82055));
	wire w61056;
	repeater #(1, 1'b0, 0, 0) c61056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61056));
	wire w69056;
	repeater #(1, 1'b0, 0, 0) c69056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69056));
	wire w77056;
	repeater #(1, 1'b0, 0, 0) c77056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77056));
	wire w58057;

	wire w59057;

	wire w63057;

	wire w66057;

	wire w67057;

	wire w71057;

	wire w74057;

	wire w75057;

	wire w79057;

	wire w58060;
	repeater #(1, 1'b0, 0, 0) c58060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58060));
	wire w63060;
	repeater #(1, 1'b0, 0, 0) c63060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63060));
	wire w74060;
	repeater #(1, 1'b0, 0, 0) c74060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74060));
	wire w79060;
	repeater #(1, 1'b0, 0, 0) c79060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79060));
	wire w58062;
	repeater #(4, 1'b0, 0, 0) c58062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58062));
	wire w63062;
	repeater #(2, 1'b0, 0, 0) c63062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63062));
	wire w64062;
	repeater #(1, 1'b0, 0, 0) c64062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64062));
	wire w66062;
	repeater #(4, 1'b0, 0, 0) c66062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66062));
	wire w74062;
	repeater #(4, 1'b0, 0, 0) c74062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74062));
	wire w79062;
	repeater #(2, 1'b0, 0, 0) c79062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79062));
	wire w66063;
	repeater #(1, 1'b0, 0, 0) c66063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66063));
	wire w70063;
	repeater #(3, 1'b0, 0, 0) c70063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70063));
	wire w63064;
	repeater #(2, 1'b0, 0, 0) c63064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63064));
	wire w79064;
	repeater #(2, 1'b0, 0, 0) c79064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79064));
	wire w71065;
	repeater #(1, 1'b0, 0, 0) c71065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71065));
	wire w72065;
	repeater #(1, 1'b0, 0, 0) c72065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72065));
	wire w61066;
	repeater #(1, 1'b0, 0, 0) c61066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61066));
	wire w69066;
	repeater #(1, 1'b0, 0, 0) c69066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69066));
	wire w71066;
	repeater #(4, 1'b0, 0, 0) c71066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71066));
	wire w77066;
	repeater #(1, 1'b0, 0, 0) c77066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77066));
	wire w58067;

	wire w59067;

	wire w63067;

	wire w66067;

	wire w67067;

	wire w71067;

	wire w74067;

	wire w75067;

	wire w79067;

	wire w91068;
	torch #(1'b1) c91068 (.i_clk(tick), .i_in(), .o_out(w91068));
	wire w58071;
	repeater #(1, 1'b0, 0, 0) c58071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58071));
	wire w59071;

	wire w62071;
	repeater #(1, 1'b0, 0, 0) c62071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62071));
	wire w63071;

	wire w66071;
	repeater #(1, 1'b0, 0, 0) c66071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66071));
	wire w67071;

	wire w70071;
	repeater #(1, 1'b0, 0, 0) c70071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70071));
	wire w71071;

	wire w74071;
	repeater #(1, 1'b0, 0, 0) c74071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74071));
	wire w75071;

	wire w78071;
	repeater #(1, 1'b0, 0, 0) c78071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78071));
	wire w79071;

	wire w82071;
	repeater #(1, 1'b0, 0, 0) c82071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82071));
	wire w83071;

	wire w58074;
	repeater #(1, 1'b0, 0, 0) c58074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58074));
	wire w63074;
	repeater #(1, 1'b0, 0, 0) c63074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63074));
	wire w66074;
	repeater #(1, 1'b0, 0, 0) c66074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66074));
	wire w71074;
	repeater #(1, 1'b0, 0, 0) c71074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71074));
	wire w74074;
	repeater #(1, 1'b0, 0, 0) c74074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74074));
	wire w79074;
	repeater #(1, 1'b0, 0, 0) c79074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79074));
	wire w82075;
	repeater #(4, 1'b0, 0, 0) c82075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82075));
	wire w58076;
	repeater #(4, 1'b0, 0, 0) c58076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58076));
	wire w63076;
	repeater #(2, 1'b0, 0, 0) c63076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63076));
	wire w66076;
	repeater #(4, 1'b0, 0, 0) c66076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66076));
	wire w71076;
	repeater #(2, 1'b0, 0, 0) c71076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71076));
	wire w74076;
	repeater #(4, 1'b0, 0, 0) c74076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74076));
	wire w79076;
	repeater #(2, 1'b0, 0, 0) c79076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79076));
	wire w63078;
	repeater #(2, 1'b0, 0, 0) c63078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63078));
	wire w71078;
	repeater #(2, 1'b0, 0, 0) c71078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71078));
	wire w79078;
	repeater #(2, 1'b0, 0, 0) c79078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79078));
	wire w82079;
	repeater #(2, 1'b0, 0, 0) c82079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82079));
	wire w61080;
	repeater #(1, 1'b0, 0, 0) c61080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61080));
	wire w69080;
	repeater #(1, 1'b0, 0, 0) c69080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69080));
	wire w77080;
	repeater #(1, 1'b0, 0, 0) c77080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77080));
	wire w58081;

	wire w59081;

	wire w63081;

	wire w66081;

	wire w67081;

	wire w71081;

	wire w74081;

	wire w75081;

	wire w79081;

	wire w58084;
	repeater #(1, 1'b0, 0, 0) c58084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58084));
	wire w63084;
	repeater #(1, 1'b0, 0, 0) c63084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63084));
	wire w74084;
	repeater #(1, 1'b0, 0, 0) c74084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74084));
	wire w79084;
	repeater #(1, 1'b0, 0, 0) c79084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79084));
	wire w58086;
	repeater #(4, 1'b0, 0, 0) c58086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58086));
	wire w63086;
	repeater #(2, 1'b0, 0, 0) c63086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63086));
	wire w64086;
	repeater #(1, 1'b0, 0, 0) c64086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w64086));
	wire w66086;
	repeater #(4, 1'b0, 0, 0) c66086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66086));
	wire w74086;
	repeater #(4, 1'b0, 0, 0) c74086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74086));
	wire w79086;
	repeater #(2, 1'b0, 0, 0) c79086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79086));
	wire w66087;
	repeater #(1, 1'b0, 0, 0) c66087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66087));
	wire w70087;
	repeater #(3, 1'b0, 0, 0) c70087 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70087));
	wire w63088;
	repeater #(2, 1'b0, 0, 0) c63088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63088));
	wire w79088;
	repeater #(2, 1'b0, 0, 0) c79088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79088));
	wire w71089;
	repeater #(1, 1'b0, 0, 0) c71089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71089));
	wire w72089;
	repeater #(1, 1'b0, 0, 0) c72089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w72089));
	wire w61090;
	repeater #(1, 1'b0, 0, 0) c61090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61090));
	wire w69090;
	repeater #(1, 1'b0, 0, 0) c69090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69090));
	wire w71090;
	repeater #(4, 1'b0, 0, 0) c71090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71090));
	wire w77090;
	repeater #(1, 1'b1, 0, 0) c77090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77090));
	wire w58091;

	wire w59091;

	wire w63091;

	wire w66091;

	wire w67091;

	wire w71091;

	wire w74091;

	wire w75091;

	wire w79091;

	wire w430145;
	repeater #(1, 1'b0, 0, 0) c430145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w430145));
	wire w540145;
	repeater #(1, 1'b0, 0, 0) c540145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540145));
	wire w540147;
	repeater #(1, 1'b0, 0, 0) c540147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540147));
	wire w580148;
	repeater #(1, 1'b0, 0, 0) c580148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580148));
	wire w380149;
	repeater #(1, 1'b0, 0, 0) c380149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380149));
	wire w390149;

	wire w570149;
	repeater #(1, 1'b0, 0, 0) c570149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w570149));
	wire w670149;
	repeater #(1, 1'b0, 0, 0) c670149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w670149));
	wire w560150;
	repeater #(1, 1'b0, 0, 0) c560150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560150));
	wire w690150;

	wire w700150;

	wire w1630150;
	repeater #(1, 1'b0, 0, 0) c1630150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630150));
	wire w1810150;
	repeater #(1, 1'b0, 0, 0) c1810150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810150));
	wire w1990150;
	repeater #(1, 1'b0, 0, 0) c1990150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990150));
	wire w90151;
	repeater #(1, 1'b0, 0, 0) c90151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90151));
	wire w270151;
	repeater #(1, 1'b0, 0, 0) c270151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w270151));
	wire w420151;

	wire w700152;
	repeater #(1, 1'b0, 0, 0) c700152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w700152));
	wire w840152;
	repeater #(1, 1'b1, 0, 0) c840152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840152));
	wire w1670152;
	repeater #(1, 1'b0, 0, 0) c1670152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1670152));
	wire w1850152;
	repeater #(1, 1'b0, 0, 0) c1850152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1850152));
	wire w2030152;
	repeater #(1, 1'b0, 0, 0) c2030152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2030152));
	wire w130153;
	repeater #(1, 1'b0, 0, 0) c130153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130153));
	wire w310153;
	repeater #(1, 1'b0, 0, 0) c310153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310153));
	wire w560153;
	repeater #(2, 1'b0, 0, 0) c560153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560153));
	wire w840153;

	wire w860154;
	repeater #(1, 1'b0, 0, 0) c860154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w860154));
	wire w560155;
	repeater #(1, 1'b0, 0, 0) c560155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560155));
	wire w900156;
	repeater #(1, 1'b1, 0, 0) c900156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w900156));
	wire w920156;
	repeater #(1, 1'b1, 0, 0) c920156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w920156));
	wire w940156;
	repeater #(1, 1'b1, 0, 0) c940156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w940156));
	wire w610162;
	repeater #(1, 1'b0, 0, 0) c610162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w610162));
	wire w690162;
	repeater #(1, 1'b0, 0, 0) c690162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w690162));
	wire w770162;
	repeater #(1, 1'b0, 0, 0) c770162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w770162));
	wire w170163;
	repeater #(1, 1'b1, 0, 0) c170163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170163));
	wire w1590164;
	repeater #(1, 1'b0, 0, 0) c1590164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1590164));
	wire w1610164;
	repeater #(1, 1'b0, 0, 0) c1610164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1610164));
	wire w860170;
	repeater #(1, 1'b0, 0, 0) c860170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w860170));
	wire w610172;
	repeater #(1, 1'b0, 0, 0) c610172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w610172));
	wire w690172;
	repeater #(1, 1'b0, 0, 0) c690172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w690172));
	wire w770172;
	repeater #(1, 1'b0, 0, 0) c770172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w770172));
	wire w900172;
	repeater #(1, 1'b1, 0, 0) c900172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w900172));
	wire w920172;
	repeater #(1, 1'b1, 0, 0) c920172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w920172));
	wire w940172;
	repeater #(1, 1'b1, 0, 0) c940172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w940172));
	wire w700176;
	repeater #(1, 1'b0, 0, 0) c700176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w700176));
	wire w840176;
	repeater #(1, 1'b1, 0, 0) c840176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w840176));
	wire w840177;

	wire w860178;
	repeater #(1, 1'b0, 0, 0) c860178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w860178));
	wire w15913;
	repeater #(1, 1'b0, 0, 0) c15913 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15913));
	wire w16113;
	repeater #(1, 1'b0, 0, 0) c16113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16113));
	wire w6117;
	repeater #(1, 1'b0, 0, 0) c6117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6117));
	wire w6917;
	repeater #(1, 1'b0, 0, 0) c6917 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6917));
	wire w7717;
	repeater #(1, 1'b0, 0, 0) c7717 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7717));
	wire w86115;
	repeater #(1, 1'b0, 0, 0) c86115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86115));
	wire w90115;
	repeater #(1, 1'b1, 0, 0) c90115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90115));
	wire w92115;
	repeater #(1, 1'b1, 0, 0) c92115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92115));
	wire w94115;
	repeater #(1, 1'b1, 0, 0) c94115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94115));
	wire w61117;
	repeater #(1, 1'b0, 0, 0) c61117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61117));
	wire w69117;
	repeater #(1, 1'b0, 0, 0) c69117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69117));
	wire w77117;
	repeater #(1, 1'b0, 0, 0) c77117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77117));
	wire w70121;
	repeater #(1, 1'b0, 0, 0) c70121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70121));
	wire w84121;
	repeater #(1, 1'b1, 0, 0) c84121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84121));
	wire w161121;
	repeater #(1, 1'b0, 0, 0) c161121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161121));
	wire w84122;

	wire w86123;
	repeater #(1, 1'b0, 0, 0) c86123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86123));
	wire w61131;
	repeater #(1, 1'b0, 0, 0) c61131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61131));
	wire w69131;
	repeater #(1, 1'b0, 0, 0) c69131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69131));
	wire w77131;
	repeater #(1, 1'b0, 0, 0) c77131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77131));
	wire w90131;
	repeater #(1, 1'b1, 0, 0) c90131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90131));
	wire w92131;
	repeater #(1, 1'b1, 0, 0) c92131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92131));
	wire w94131;
	repeater #(1, 1'b1, 0, 0) c94131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94131));
	wire w86139;
	repeater #(1, 1'b0, 0, 0) c86139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86139));
	wire w61141;
	repeater #(1, 1'b0, 0, 0) c61141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61141));
	wire w69141;
	repeater #(1, 1'b0, 0, 0) c69141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69141));
	wire w77141;
	repeater #(1, 1'b0, 0, 0) c77141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77141));
	wire w70145;
	repeater #(1, 1'b0, 0, 0) c70145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70145));
	wire w84145;
	repeater #(1, 1'b1, 0, 0) c84145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84145));
	wire w84146;

	wire w86147;
	repeater #(1, 1'b0, 0, 0) c86147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86147));
	wire w90147;
	repeater #(1, 1'b1, 0, 0) c90147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90147));
	wire w92147;
	repeater #(1, 1'b1, 0, 0) c92147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92147));
	wire w94147;
	repeater #(1, 1'b1, 0, 0) c94147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94147));
	wire w61155;
	repeater #(1, 1'b0, 0, 0) c61155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61155));
	wire w69155;
	repeater #(1, 1'b0, 0, 0) c69155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69155));
	wire w77155;
	repeater #(1, 1'b0, 0, 0) c77155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77155));
	wire w86163;
	repeater #(1, 1'b0, 0, 0) c86163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86163));
	wire w90163;
	repeater #(1, 1'b1, 0, 0) c90163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90163));
	wire w92163;
	repeater #(1, 1'b1, 0, 0) c92163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w92163));
	wire w94163;
	repeater #(1, 1'b1, 0, 0) c94163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94163));
	wire w61165;
	repeater #(1, 1'b0, 0, 0) c61165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61165));
	wire w69165;
	repeater #(1, 1'b0, 0, 0) c69165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69165));
	wire w77165;
	repeater #(1, 1'b0, 0, 0) c77165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77165));
	wire w70169;
	repeater #(1, 1'b0, 0, 0) c70169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70169));
	wire w84169;
	repeater #(1, 1'b1, 0, 0) c84169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w84169));
	wire w84170;

	wire w86171;
	repeater #(1, 1'b0, 0, 0) c86171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86171));
	wire w61179;
	repeater #(1, 1'b0, 0, 0) c61179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61179));
	wire w69179;
	repeater #(1, 1'b0, 0, 0) c69179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69179));
	wire w77179;
	repeater #(1, 1'b0, 0, 0) c77179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77179));
	wire w86187;
	repeater #(1, 1'b0, 0, 0) c86187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86187));
	wire w61189;
	repeater #(1, 1'b0, 0, 0) c61189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w61189));
	wire w69189;
	repeater #(1, 1'b0, 0, 0) c69189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w69189));
	wire w77189;
	repeater #(1, 1'b0, 0, 0) c77189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w77189));
	wire w88192;
	repeater #(1, 1'b0, 0, 0) c88192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w88192));
	wire w70193;
	repeater #(1, 1'b0, 0, 0) c70193 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70193));
	wire w89194;

	wire w92194;
	assign outputs[118] = ();
	wire w89195;

	wire w87196;
	repeater #(1, 1'b0, 0, 0) c87196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87196));
	wire w58198;
	repeater #(1, 1'b0, 0, 0) c58198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58198));
	wire w62198;
	repeater #(1, 1'b0, 0, 0) c62198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62198));
	wire w66198;
	repeater #(1, 1'b0, 0, 0) c66198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66198));
	wire w70198;
	repeater #(1, 1'b0, 0, 0) c70198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70198));
	wire w74198;
	repeater #(1, 1'b0, 0, 0) c74198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74198));
	wire w78198;
	repeater #(1, 1'b0, 0, 0) c78198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78198));
	wire w82198;
	repeater #(1, 1'b0, 0, 0) c82198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82198));
	wire w33016;
	repeater #(1, 1'b0, 0, 0) c33016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33016));
	wire w42018;
	repeater #(1, 1'b1, 0, 0) c42018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42018));
	wire w43018;

	wire w46018;
	repeater #(1, 1'b1, 0, 0) c46018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46018));
	wire w47018;

	wire w50018;
	repeater #(1, 1'b1, 0, 0) c50018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50018));
	wire w51018;

	wire w54018;
	repeater #(1, 1'b1, 0, 0) c54018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54018));
	wire w55018;

	wire w58018;
	repeater #(1, 1'b1, 0, 0) c58018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58018));
	wire w59018;

	wire w62018;
	repeater #(1, 1'b0, 0, 0) c62018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62018));
	wire w63018;

	wire w66018;
	repeater #(1, 1'b1, 0, 0) c66018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66018));
	wire w67018;

	wire w33019;
	repeater #(2, 1'b0, 0, 0) c33019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33019));
	wire w35019;
	repeater #(2, 1'b0, 0, 0) c35019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35019));
	wire w37019;
	repeater #(2, 1'b0, 0, 0) c37019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37019));
	wire w35020;
	repeater #(2, 1'b0, 0, 0) c35020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35020));
	wire w37020;
	repeater #(2, 1'b0, 0, 0) c37020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37020));
	wire w35021;
	repeater #(2, 1'b0, 0, 0) c35021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35021));
	wire w37021;
	repeater #(2, 1'b0, 0, 0) c37021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37021));
	wire w42021;
	repeater #(1, 1'b1, 0, 0) c42021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42021));
	wire w47021;
	repeater #(1, 1'b1, 0, 0) c47021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47021));
	wire w50021;
	repeater #(1, 1'b1, 0, 0) c50021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50021));
	wire w55021;
	repeater #(1, 1'b1, 0, 0) c55021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55021));
	wire w58021;
	repeater #(1, 1'b1, 0, 0) c58021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58021));
	wire w63021;
	repeater #(1, 1'b0, 0, 0) c63021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63021));
	wire w35022;
	repeater #(2, 1'b0, 0, 0) c35022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35022));
	wire w37022;
	repeater #(2, 1'b0, 0, 0) c37022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37022));
	wire w39022;
	repeater #(1, 1'b0, 0, 0) c39022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39022));
	wire w44022;

	wire w45022;

	wire w52022;

	wire w53022;

	wire w60022;

	wire w61022;

	wire w66022;
	repeater #(4, 1'b1, 0, 0) c66022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66022));
	wire w35023;
	repeater #(1, 1'b0, 0, 0) c35023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35023));
	wire w37023;
	repeater #(1, 1'b0, 0, 0) c37023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37023));
	wire w39023;
	repeater #(1, 1'b0, 0, 0) c39023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39023));
	wire w42023;
	repeater #(4, 1'b1, 0, 0) c42023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42023));
	wire w47023;
	repeater #(2, 1'b1, 0, 0) c47023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47023));
	wire w50023;
	repeater #(4, 1'b1, 0, 0) c50023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50023));
	wire w55023;
	repeater #(2, 1'b1, 0, 0) c55023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55023));
	wire w58023;
	repeater #(4, 1'b1, 0, 0) c58023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58023));
	wire w63023;
	repeater #(2, 1'b0, 0, 0) c63023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63023));
	wire w33024;
	repeater #(2, 1'b0, 0, 0) c33024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33024));
	wire w39024;
	repeater #(2, 1'b0, 0, 0) c39024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39024));
	wire w35025;
	repeater #(1, 1'b0, 0, 0) c35025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35025));
	wire w37025;
	repeater #(1, 1'b0, 0, 0) c37025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37025));
	wire w47025;
	repeater #(2, 1'b1, 0, 0) c47025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47025));
	wire w55025;
	repeater #(2, 1'b1, 0, 0) c55025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55025));
	wire w63025;
	repeater #(2, 1'b0, 0, 0) c63025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63025));
	wire w2026;

	wire w66026;
	repeater #(2, 1'b1, 0, 0) c66026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66026));
	wire w42028;

	wire w43028;

	wire w46028;
	repeater #(1, 1'b0, 0, 0) c46028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46028));
	wire w47028;

	wire w50028;

	wire w51028;

	wire w54028;
	repeater #(1, 1'b1, 0, 0) c54028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54028));
	wire w55028;

	wire w58028;

	wire w59028;

	wire w62028;
	repeater #(1, 1'b1, 0, 0) c62028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62028));
	wire w63028;

	wire w42031;
	repeater #(1, 1'b1, 0, 0) c42031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42031));
	wire w47031;
	repeater #(1, 1'b1, 0, 0) c47031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47031));
	wire w58031;
	repeater #(1, 1'b1, 0, 0) c58031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58031));
	wire w63031;
	repeater #(1, 1'b1, 0, 0) c63031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63031));
	wire w44032;

	wire w45032;

	wire w49032;
	repeater #(1, 1'b1, 0, 0) c49032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49032));
	wire w52032;

	wire w53032;

	wire w60032;

	wire w61032;

	wire w42033;
	repeater #(4, 1'b1, 0, 0) c42033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42033));
	wire w47033;
	repeater #(2, 1'b1, 0, 0) c47033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47033));
	wire w48033;
	repeater #(1, 1'b1, 0, 0) c48033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48033));
	wire w50033;
	repeater #(4, 1'b1, 0, 0) c50033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50033));
	wire w55033;
	repeater #(1, 1'b1, 0, 0) c55033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55033));
	wire w58033;
	repeater #(4, 1'b1, 0, 0) c58033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58033));
	wire w63033;
	repeater #(2, 1'b1, 0, 0) c63033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63033));
	wire w47035;
	repeater #(2, 1'b1, 0, 0) c47035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47035));
	wire w63035;
	repeater #(2, 1'b1, 0, 0) c63035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63035));
	wire w55036;
	repeater #(1, 1'b1, 0, 0) c55036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55036));
	wire w56036;
	repeater #(1, 1'b1, 0, 0) c56036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56036));
	wire w55037;
	repeater #(4, 1'b1, 0, 0) c55037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55037));
	wire w42038;

	wire w43038;

	wire w46038;
	repeater #(1, 1'b0, 0, 0) c46038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46038));
	wire w47038;

	wire w50038;

	wire w51038;

	wire w54038;
	repeater #(1, 1'b1, 0, 0) c54038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54038));
	wire w55038;

	wire w58038;

	wire w59038;

	wire w62038;
	repeater #(1, 1'b1, 0, 0) c62038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62038));
	wire w63038;

	wire w56040;
	torch #(1'b1) c56040 (.i_clk(tick), .i_in(), .o_out(w56040));
	wire w42042;
	repeater #(1, 1'b1, 0, 0) c42042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42042));
	wire w43042;

	wire w46042;
	repeater #(1, 1'b0, 0, 0) c46042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46042));
	wire w47042;

	wire w50042;
	repeater #(1, 1'b0, 0, 0) c50042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50042));
	wire w51042;

	wire w54042;
	repeater #(1, 1'b1, 0, 0) c54042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54042));
	wire w55042;

	wire w58042;
	repeater #(1, 1'b0, 0, 0) c58042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58042));
	wire w59042;

	wire w62042;
	repeater #(1, 1'b0, 0, 0) c62042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62042));
	wire w63042;

	wire w66042;
	repeater #(1, 1'b0, 0, 0) c66042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66042));
	wire w67042;

	wire w42045;
	repeater #(1, 1'b1, 0, 0) c42045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42045));
	wire w47045;
	repeater #(1, 1'b0, 0, 0) c47045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47045));
	wire w50045;
	repeater #(1, 1'b0, 0, 0) c50045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50045));
	wire w55045;
	repeater #(1, 1'b1, 0, 0) c55045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55045));
	wire w58045;
	repeater #(1, 1'b0, 0, 0) c58045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58045));
	wire w63045;
	repeater #(1, 1'b0, 0, 0) c63045 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63045));
	wire w44046;

	wire w45046;

	wire w52046;

	wire w53046;

	wire w60046;

	wire w61046;

	wire w66046;
	repeater #(4, 1'b0, 0, 0) c66046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66046));
	wire w42047;
	repeater #(4, 1'b1, 0, 0) c42047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42047));
	wire w47047;
	repeater #(2, 1'b0, 0, 0) c47047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47047));
	wire w50047;
	repeater #(4, 1'b0, 0, 0) c50047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50047));
	wire w55047;
	repeater #(2, 1'b1, 0, 0) c55047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55047));
	wire w58047;
	repeater #(4, 1'b0, 0, 0) c58047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58047));
	wire w63047;
	repeater #(2, 1'b0, 0, 0) c63047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63047));
	wire w47049;
	repeater #(2, 1'b0, 0, 0) c47049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47049));
	wire w55049;
	repeater #(2, 1'b1, 0, 0) c55049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55049));
	wire w63049;
	repeater #(2, 1'b0, 0, 0) c63049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63049));
	wire w66050;
	repeater #(2, 1'b0, 0, 0) c66050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66050));
	wire w42052;

	wire w43052;

	wire w46052;
	repeater #(1, 1'b1, 0, 0) c46052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46052));
	wire w47052;

	wire w50052;

	wire w51052;

	wire w54052;
	repeater #(1, 1'b0, 0, 0) c54052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54052));
	wire w55052;

	wire w58052;

	wire w59052;

	wire w62052;
	repeater #(1, 1'b1, 0, 0) c62052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62052));
	wire w63052;

	wire w42055;
	repeater #(1, 1'b1, 0, 0) c42055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42055));
	wire w47055;
	repeater #(1, 1'b1, 0, 0) c47055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47055));
	wire w58055;
	repeater #(1, 1'b0, 0, 0) c58055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58055));
	wire w63055;
	repeater #(1, 1'b0, 0, 0) c63055 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63055));
	wire w44056;

	wire w45056;

	wire w49056;
	repeater #(1, 1'b1, 0, 0) c49056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49056));
	wire w52056;

	wire w53056;

	wire w60056;

	wire w61056;

	wire w42057;
	repeater #(4, 1'b1, 0, 0) c42057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42057));
	wire w47057;
	repeater #(2, 1'b1, 0, 0) c47057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47057));
	wire w48057;
	repeater #(1, 1'b1, 0, 0) c48057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48057));
	wire w50057;
	repeater #(4, 1'b1, 0, 0) c50057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50057));
	wire w55057;
	repeater #(1, 1'b0, 0, 0) c55057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55057));
	wire w58057;
	repeater #(4, 1'b0, 0, 0) c58057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58057));
	wire w63057;
	repeater #(2, 1'b0, 0, 0) c63057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63057));
	wire w47059;
	repeater #(2, 1'b1, 0, 0) c47059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47059));
	wire w63059;
	repeater #(2, 1'b0, 0, 0) c63059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63059));
	wire w55060;
	repeater #(1, 1'b0, 0, 0) c55060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55060));
	wire w56060;
	repeater #(1, 1'b0, 0, 0) c56060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56060));
	wire w55061;
	repeater #(4, 1'b0, 0, 0) c55061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55061));
	wire w42062;

	wire w43062;

	wire w46062;
	repeater #(1, 1'b0, 0, 0) c46062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46062));
	wire w47062;

	wire w50062;

	wire w51062;

	wire w54062;
	repeater #(1, 1'b1, 0, 0) c54062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54062));
	wire w55062;

	wire w58062;

	wire w59062;

	wire w62062;
	repeater #(1, 1'b1, 0, 0) c62062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62062));
	wire w63062;

	wire w56064;
	torch #(1'b1) c56064 (.i_clk(tick), .i_in(), .o_out(w56064));
	wire w42066;
	repeater #(1, 1'b0, 0, 0) c42066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42066));
	wire w43066;

	wire w46066;
	repeater #(1, 1'b0, 0, 0) c46066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46066));
	wire w47066;

	wire w50066;
	repeater #(1, 1'b0, 0, 0) c50066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50066));
	wire w51066;

	wire w54066;
	repeater #(1, 1'b0, 0, 0) c54066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54066));
	wire w55066;

	wire w58066;
	repeater #(1, 1'b0, 0, 0) c58066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58066));
	wire w59066;

	wire w62066;
	repeater #(1, 1'b1, 0, 0) c62066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62066));
	wire w63066;

	wire w66066;
	repeater #(1, 1'b0, 0, 0) c66066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66066));
	wire w67066;

	wire w42069;
	repeater #(1, 1'b0, 0, 0) c42069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42069));
	wire w47069;
	repeater #(1, 1'b0, 0, 0) c47069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47069));
	wire w50069;
	repeater #(1, 1'b0, 0, 0) c50069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50069));
	wire w55069;
	repeater #(1, 1'b0, 0, 0) c55069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55069));
	wire w58069;
	repeater #(1, 1'b0, 0, 0) c58069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58069));
	wire w63069;
	repeater #(1, 1'b1, 0, 0) c63069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63069));
	wire w44070;

	wire w45070;

	wire w52070;

	wire w53070;

	wire w60070;

	wire w61070;

	wire w66070;
	repeater #(4, 1'b0, 0, 0) c66070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66070));
	wire w42071;
	repeater #(4, 1'b0, 0, 0) c42071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42071));
	wire w47071;
	repeater #(2, 1'b0, 0, 0) c47071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47071));
	wire w50071;
	repeater #(4, 1'b0, 0, 0) c50071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50071));
	wire w55071;
	repeater #(2, 1'b0, 0, 0) c55071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55071));
	wire w58071;
	repeater #(4, 1'b0, 0, 0) c58071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58071));
	wire w63071;
	repeater #(2, 1'b1, 0, 0) c63071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63071));
	wire w47073;
	repeater #(2, 1'b0, 0, 0) c47073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47073));
	wire w55073;
	repeater #(2, 1'b0, 0, 0) c55073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55073));
	wire w63073;
	repeater #(2, 1'b1, 0, 0) c63073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63073));
	wire w66074;
	repeater #(2, 1'b0, 0, 0) c66074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66074));
	wire w42076;

	wire w43076;

	wire w46076;
	repeater #(1, 1'b0, 0, 0) c46076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46076));
	wire w47076;

	wire w50076;

	wire w51076;

	wire w54076;
	repeater #(1, 1'b0, 0, 0) c54076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54076));
	wire w55076;

	wire w58076;

	wire w59076;

	wire w62076;
	repeater #(1, 1'b1, 0, 0) c62076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62076));
	wire w63076;

	wire w42079;
	repeater #(1, 1'b0, 0, 0) c42079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42079));
	wire w47079;
	repeater #(1, 1'b0, 0, 0) c47079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47079));
	wire w58079;
	repeater #(1, 1'b0, 0, 0) c58079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58079));
	wire w63079;
	repeater #(1, 1'b0, 0, 0) c63079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63079));
	wire w44080;

	wire w45080;

	wire w49080;
	repeater #(1, 1'b0, 0, 0) c49080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w49080));
	wire w52080;

	wire w53080;

	wire w60080;

	wire w61080;

	wire w42081;
	repeater #(4, 1'b0, 0, 0) c42081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42081));
	wire w47081;
	repeater #(2, 1'b0, 0, 0) c47081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47081));
	wire w48081;
	repeater #(1, 1'b0, 0, 0) c48081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w48081));
	wire w50081;
	repeater #(4, 1'b0, 0, 0) c50081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50081));
	wire w55081;
	repeater #(1, 1'b0, 0, 0) c55081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55081));
	wire w58081;
	repeater #(4, 1'b0, 0, 0) c58081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58081));
	wire w63081;
	repeater #(2, 1'b0, 0, 0) c63081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63081));
	wire w47083;
	repeater #(2, 1'b0, 0, 0) c47083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47083));
	wire w63083;
	repeater #(2, 1'b0, 0, 0) c63083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63083));
	wire w55084;
	repeater #(1, 1'b0, 0, 0) c55084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55084));
	wire w56084;
	repeater #(1, 1'b0, 0, 0) c56084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56084));
	wire w55085;
	repeater #(4, 1'b0, 0, 0) c55085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55085));
	wire w42086;

	wire w43086;

	wire w46086;
	repeater #(1, 1'b0, 0, 0) c46086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46086));
	wire w47086;

	wire w50086;

	wire w51086;

	wire w54086;
	repeater #(1, 1'b1, 0, 0) c54086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54086));
	wire w55086;

	wire w58086;

	wire w59086;

	wire w62086;
	repeater #(1, 1'b1, 0, 0) c62086 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62086));
	wire w63086;

	wire w56088;
	torch #(1'b0) c56088 (.i_clk(tick), .i_in(), .o_out(w56088));
	wire w42090;
	repeater #(1, 1'b0, 0, 0) c42090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42090));
	wire w43090;

	wire w46090;
	repeater #(1, 1'b0, 0, 0) c46090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46090));
	wire w47090;

	wire w50090;
	repeater #(1, 1'b0, 0, 0) c50090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50090));
	wire w51090;

	wire w54090;
	repeater #(1, 1'b0, 0, 0) c54090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54090));
	wire w55090;

	wire w58090;
	repeater #(1, 1'b0, 0, 0) c58090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58090));
	wire w59090;

	wire w62090;
	repeater #(1, 1'b0, 0, 0) c62090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w62090));
	wire w63090;

	wire w66090;
	repeater #(1, 1'b0, 0, 0) c66090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66090));
	wire w67090;

	wire w42093;
	repeater #(1, 1'b0, 0, 0) c42093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42093));
	wire w47093;
	repeater #(1, 1'b0, 0, 0) c47093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47093));
	wire w50093;
	repeater #(1, 1'b0, 0, 0) c50093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50093));
	wire w55093;
	repeater #(1, 1'b0, 0, 0) c55093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55093));
	wire w58093;
	repeater #(1, 1'b0, 0, 0) c58093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58093));
	wire w63093;
	repeater #(1, 1'b0, 0, 0) c63093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63093));
	wire w44094;

	wire w45094;

	wire w52094;

	wire w53094;

	wire w60094;

	wire w61094;

	wire w66094;
	repeater #(4, 1'b0, 0, 0) c66094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66094));
	wire w42095;
	repeater #(4, 1'b0, 0, 0) c42095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42095));
	wire w47095;
	repeater #(2, 1'b0, 0, 0) c47095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47095));
	wire w50095;
	repeater #(4, 1'b0, 0, 0) c50095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50095));
	wire w55095;
	repeater #(2, 1'b0, 0, 0) c55095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55095));
	wire w58095;
	repeater #(4, 1'b0, 0, 0) c58095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w58095));
	wire w63095;
	repeater #(2, 1'b0, 0, 0) c63095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63095));
	wire w47097;
	repeater #(2, 1'b0, 0, 0) c47097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47097));
	wire w55097;
	repeater #(2, 1'b0, 0, 0) c55097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w55097));
	wire w63097;
	repeater #(2, 1'b0, 0, 0) c63097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w63097));
	wire w66098;
	repeater #(2, 1'b0, 0, 0) c66098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w66098));
	wire w420100;

	wire w430100;

	wire w460100;
	repeater #(1, 1'b0, 0, 0) c460100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460100));
	wire w470100;

	wire w500100;

	wire w510100;

	wire w540100;
	repeater #(1, 1'b0, 0, 0) c540100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540100));
	wire w550100;

	wire w580100;

	wire w590100;

	wire w620100;
	repeater #(1, 1'b0, 0, 0) c620100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620100));
	wire w630100;

	wire w420103;
	repeater #(1, 1'b0, 0, 0) c420103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420103));
	wire w470103;
	repeater #(1, 1'b0, 0, 0) c470103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470103));
	wire w580103;
	repeater #(1, 1'b0, 0, 0) c580103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580103));
	wire w630103;
	repeater #(1, 1'b0, 0, 0) c630103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630103));
	wire w440104;

	wire w450104;

	wire w490104;
	repeater #(1, 1'b0, 0, 0) c490104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w490104));
	wire w520104;

	wire w530104;

	wire w600104;

	wire w610104;

	wire w420105;
	repeater #(4, 1'b0, 0, 0) c420105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420105));
	wire w470105;
	repeater #(2, 1'b0, 0, 0) c470105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470105));
	wire w480105;
	repeater #(1, 1'b0, 0, 0) c480105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480105));
	wire w500105;
	repeater #(4, 1'b0, 0, 0) c500105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500105));
	wire w550105;
	repeater #(1, 1'b0, 0, 0) c550105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550105));
	wire w580105;
	repeater #(4, 1'b0, 0, 0) c580105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580105));
	wire w630105;
	repeater #(2, 1'b0, 0, 0) c630105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630105));
	wire w470107;
	repeater #(2, 1'b0, 0, 0) c470107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470107));
	wire w630107;
	repeater #(2, 1'b0, 0, 0) c630107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630107));
	wire w550108;
	repeater #(1, 1'b0, 0, 0) c550108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550108));
	wire w560108;
	repeater #(1, 1'b0, 0, 0) c560108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560108));
	wire w550109;
	repeater #(4, 1'b0, 0, 0) c550109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550109));
	wire w420110;

	wire w430110;

	wire w460110;
	repeater #(1, 1'b0, 0, 0) c460110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460110));
	wire w470110;

	wire w500110;

	wire w510110;

	wire w540110;
	repeater #(1, 1'b0, 0, 0) c540110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540110));
	wire w550110;

	wire w580110;

	wire w590110;

	wire w620110;
	repeater #(1, 1'b0, 0, 0) c620110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620110));
	wire w630110;

	wire w560112;
	torch #(1'b0) c560112 (.i_clk(tick), .i_in(), .o_out(w560112));
	wire w420114;
	repeater #(1, 1'b1, 0, 0) c420114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420114));
	wire w430114;

	wire w460114;
	repeater #(1, 1'b1, 0, 0) c460114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460114));
	wire w470114;

	wire w500114;
	repeater #(1, 1'b1, 0, 0) c500114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500114));
	wire w510114;

	wire w540114;
	repeater #(1, 1'b1, 0, 0) c540114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540114));
	wire w550114;

	wire w580114;
	repeater #(1, 1'b1, 0, 0) c580114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580114));
	wire w590114;

	wire w620114;
	repeater #(1, 1'b1, 0, 0) c620114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620114));
	wire w630114;

	wire w660114;
	repeater #(1, 1'b1, 0, 0) c660114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660114));
	wire w670114;

	wire w420117;
	repeater #(1, 1'b1, 0, 0) c420117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420117));
	wire w470117;
	repeater #(1, 1'b1, 0, 0) c470117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470117));
	wire w500117;
	repeater #(1, 1'b1, 0, 0) c500117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500117));
	wire w550117;
	repeater #(1, 1'b1, 0, 0) c550117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550117));
	wire w580117;
	repeater #(1, 1'b1, 0, 0) c580117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580117));
	wire w630117;
	repeater #(1, 1'b1, 0, 0) c630117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630117));
	wire w440118;

	wire w450118;

	wire w520118;

	wire w530118;

	wire w600118;

	wire w610118;

	wire w660118;
	repeater #(4, 1'b1, 0, 0) c660118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660118));
	wire w420119;
	repeater #(4, 1'b1, 0, 0) c420119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420119));
	wire w470119;
	repeater #(2, 1'b1, 0, 0) c470119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470119));
	wire w500119;
	repeater #(4, 1'b1, 0, 0) c500119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500119));
	wire w550119;
	repeater #(2, 1'b1, 0, 0) c550119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550119));
	wire w580119;
	repeater #(4, 1'b1, 0, 0) c580119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580119));
	wire w630119;
	repeater #(2, 1'b1, 0, 0) c630119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630119));
	wire w470121;
	repeater #(2, 1'b1, 0, 0) c470121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470121));
	wire w550121;
	repeater #(2, 1'b1, 0, 0) c550121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550121));
	wire w630121;
	repeater #(2, 1'b1, 0, 0) c630121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630121));
	wire w660122;
	repeater #(2, 1'b1, 0, 0) c660122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w660122));
	wire w420124;

	wire w430124;

	wire w460124;
	repeater #(1, 1'b0, 0, 0) c460124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460124));
	wire w470124;

	wire w500124;

	wire w510124;

	wire w540124;
	repeater #(1, 1'b0, 0, 0) c540124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540124));
	wire w550124;

	wire w580124;

	wire w590124;

	wire w620124;
	repeater #(1, 1'b0, 0, 0) c620124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620124));
	wire w630124;

	wire w420127;
	repeater #(1, 1'b1, 0, 0) c420127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420127));
	wire w470127;
	repeater #(1, 1'b1, 0, 0) c470127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470127));
	wire w580127;
	repeater #(1, 1'b1, 0, 0) c580127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580127));
	wire w630127;
	repeater #(1, 1'b1, 0, 0) c630127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630127));
	wire w440128;

	wire w450128;

	wire w490128;
	repeater #(1, 1'b1, 0, 0) c490128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w490128));
	wire w520128;

	wire w530128;

	wire w600128;

	wire w610128;

	wire w420129;
	repeater #(4, 1'b1, 0, 0) c420129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420129));
	wire w470129;
	repeater #(2, 1'b1, 0, 0) c470129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470129));
	wire w480129;
	repeater #(1, 1'b1, 0, 0) c480129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w480129));
	wire w500129;
	repeater #(4, 1'b1, 0, 0) c500129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500129));
	wire w550129;
	repeater #(1, 1'b1, 0, 0) c550129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550129));
	wire w580129;
	repeater #(4, 1'b1, 0, 0) c580129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w580129));
	wire w630129;
	repeater #(2, 1'b1, 0, 0) c630129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630129));
	wire w470131;
	repeater #(2, 1'b1, 0, 0) c470131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470131));
	wire w630131;
	repeater #(2, 1'b1, 0, 0) c630131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w630131));
	wire w550132;
	repeater #(1, 1'b1, 0, 0) c550132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550132));
	wire w560132;
	repeater #(1, 1'b1, 0, 0) c560132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w560132));
	wire w550133;
	repeater #(4, 1'b1, 0, 0) c550133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w550133));
	wire w420134;

	wire w430134;

	wire w460134;
	repeater #(1, 1'b0, 0, 0) c460134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460134));
	wire w470134;

	wire w500134;

	wire w510134;

	wire w540134;
	repeater #(1, 1'b0, 0, 0) c540134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w540134));
	wire w550134;

	wire w580134;

	wire w590134;

	wire w620134;
	repeater #(1, 1'b1, 0, 0) c620134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w620134));
	wire w630134;

	wire w560136;
	torch #(1'b1) c560136 (.i_clk(tick), .i_in(), .o_out(w560136));
	wire w41111;
	repeater #(1, 1'b0, 0, 0) c41111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41111));
	wire w42112;
	repeater #(1, 1'b0, 0, 0) c42112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42112));
	wire w4113;
	repeater #(1, 1'b1, 0, 0) c4113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4113));
	wire w21113;
	repeater #(2, 1'b1, 0, 0) c21113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21113));
	wire w22113;
	repeater #(1, 1'b1, 0, 0) c22113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22113));
	wire w23113;

	wire w38113;

	wire w41113;
	repeater #(1, 1'b1, 0, 0) c41113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w41113));
	wire w51113;
	repeater #(1, 1'b1, 0, 0) c51113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w51113));
	wire w56113;
	repeater #(1, 1'b1, 0, 0) c56113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w56113));
	wire w40114;
	repeater #(1, 1'b0, 0, 0) c40114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40114));
	wire w53114;

	wire w54114;

	wire w37115;
	repeater #(1, 1'b0, 0, 0) c37115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w37115));
	wire w54116;
	repeater #(1, 1'b0, 0, 0) c54116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54116));
	wire w68116;
	repeater #(1, 1'b1, 0, 0) c68116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68116));
	wire w68117;

	wire w70118;
	repeater #(1, 1'b0, 0, 0) c70118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70118));
	wire w39119;
	repeater #(1, 1'b0, 0, 0) c39119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39119));
	wire w2127;
	repeater #(1, 1'b0, 0, 0) c2127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2127));
	wire w70134;
	repeater #(1, 1'b0, 0, 0) c70134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70134));
	wire w68140;
	repeater #(1, 1'b1, 0, 0) c68140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68140));
	wire w68141;

	wire w70142;
	repeater #(1, 1'b0, 0, 0) c70142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70142));
	wire w70158;
	repeater #(1, 1'b0, 0, 0) c70158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70158));
	wire w68164;
	repeater #(1, 1'b1, 0, 0) c68164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68164));
	wire w68165;

	wire w70166;
	repeater #(1, 1'b0, 0, 0) c70166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70166));
	wire w70182;
	repeater #(1, 1'b0, 0, 0) c70182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70182));
	wire w68188;
	repeater #(1, 1'b1, 0, 0) c68188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w68188));
	wire w68189;

	wire w70190;
	repeater #(1, 1'b0, 0, 0) c70190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70190));
	wire w701106;
	repeater #(1, 1'b0, 0, 0) c701106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w701106));
	wire w681112;
	repeater #(1, 1'b1, 0, 0) c681112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w681112));
	wire w681113;

	wire w701114;
	repeater #(1, 1'b0, 0, 0) c701114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w701114));
	wire w701130;
	repeater #(1, 1'b0, 0, 0) c701130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w701130));
	wire w721135;
	repeater #(1, 1'b0, 0, 0) c721135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w721135));
	wire w5701;

	wire w6001;
	assign outputs[119] = ();
	wire w5702;

	wire w5503;
	repeater #(1, 1'b0, 0, 0) c5503 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5503));
	wire w197055;

	wire w20060;
	repeater #(1, 1'b0, 0, 0) c20060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20060));
	wire w26061;
	repeater #(1, 1'b1, 0, 0) c26061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26061));
	wire w27061;

	wire w30061;
	repeater #(1, 1'b0, 0, 0) c30061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30061));
	wire w31061;

	wire w34061;
	repeater #(1, 1'b0, 0, 0) c34061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34061));
	wire w35061;

	wire w38061;
	repeater #(1, 1'b1, 0, 0) c38061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38061));
	wire w39061;

	wire w42061;
	repeater #(1, 1'b1, 0, 0) c42061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42061));
	wire w43061;

	wire w46061;
	repeater #(1, 1'b1, 0, 0) c46061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46061));
	wire w47061;

	wire w50061;
	repeater #(1, 1'b0, 0, 0) c50061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50061));
	wire w51061;

	wire w19062;
	repeater #(2, 1'b0, 0, 0) c19062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19062));
	wire w21063;
	repeater #(1, 1'b0, 0, 0) c21063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21063));
	wire w19064;
	repeater #(2, 1'b0, 0, 0) c19064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19064));
	wire w21064;
	repeater #(2, 1'b0, 0, 0) c21064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21064));
	wire w26064;
	repeater #(1, 1'b1, 0, 0) c26064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26064));
	wire w31064;
	repeater #(1, 1'b0, 0, 0) c31064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31064));
	wire w34064;
	repeater #(1, 1'b0, 0, 0) c34064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34064));
	wire w39064;
	repeater #(1, 1'b1, 0, 0) c39064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39064));
	wire w42064;
	repeater #(1, 1'b1, 0, 0) c42064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42064));
	wire w47064;
	repeater #(1, 1'b1, 0, 0) c47064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47064));
	wire w21065;
	repeater #(2, 1'b0, 0, 0) c21065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21065));
	wire w28065;

	wire w29065;

	wire w36065;

	wire w37065;

	wire w44065;

	wire w45065;

	wire w50065;
	repeater #(4, 1'b0, 0, 0) c50065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50065));
	wire w26066;
	repeater #(4, 1'b1, 0, 0) c26066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26066));
	wire w31066;
	repeater #(2, 1'b0, 0, 0) c31066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31066));
	wire w34066;
	repeater #(4, 1'b0, 0, 0) c34066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34066));
	wire w39066;
	repeater #(2, 1'b1, 0, 0) c39066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39066));
	wire w42066;
	repeater #(4, 1'b1, 0, 0) c42066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42066));
	wire w47066;
	repeater #(2, 1'b1, 0, 0) c47066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47066));
	wire w31068;
	repeater #(2, 1'b0, 0, 0) c31068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31068));
	wire w39068;
	repeater #(2, 1'b1, 0, 0) c39068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39068));
	wire w47068;
	repeater #(2, 1'b1, 0, 0) c47068 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47068));
	wire w193068;

	wire w50069;
	repeater #(2, 1'b0, 0, 0) c50069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50069));
	wire w26071;

	wire w27071;

	wire w30071;
	repeater #(1, 1'b0, 0, 0) c30071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30071));
	wire w31071;

	wire w34071;

	wire w35071;

	wire w38071;
	repeater #(1, 1'b1, 0, 0) c38071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38071));
	wire w39071;

	wire w42071;

	wire w43071;

	wire w46071;
	repeater #(1, 1'b1, 0, 0) c46071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46071));
	wire w47071;

	wire w26074;
	repeater #(1, 1'b0, 0, 0) c26074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26074));
	wire w31074;
	repeater #(1, 1'b0, 0, 0) c31074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31074));
	wire w42074;
	repeater #(1, 1'b1, 0, 0) c42074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42074));
	wire w47074;
	repeater #(1, 1'b0, 0, 0) c47074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47074));
	wire w28075;

	wire w29075;

	wire w33075;
	repeater #(1, 1'b0, 0, 0) c33075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33075));
	wire w36075;

	wire w37075;

	wire w44075;

	wire w45075;

	wire w26076;
	repeater #(4, 1'b0, 0, 0) c26076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26076));
	wire w31076;
	repeater #(2, 1'b0, 0, 0) c31076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31076));
	wire w32076;
	repeater #(1, 1'b0, 0, 0) c32076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w32076));
	wire w34076;
	repeater #(4, 1'b0, 0, 0) c34076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34076));
	wire w39076;
	repeater #(1, 1'b1, 0, 0) c39076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39076));
	wire w42076;
	repeater #(4, 1'b1, 0, 0) c42076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42076));
	wire w47076;
	repeater #(2, 1'b0, 0, 0) c47076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47076));
	wire w31078;
	repeater #(2, 1'b0, 0, 0) c31078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31078));
	wire w47078;
	repeater #(2, 1'b0, 0, 0) c47078 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47078));
	wire w39079;
	repeater #(1, 1'b1, 0, 0) c39079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39079));
	wire w40079;
	repeater #(1, 1'b1, 0, 0) c40079 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40079));
	wire w39080;
	repeater #(4, 1'b1, 0, 0) c39080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39080));
	wire w26081;

	wire w27081;

	wire w30081;
	repeater #(1, 1'b0, 0, 0) c30081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30081));
	wire w31081;

	wire w34081;

	wire w35081;

	wire w38081;
	repeater #(1, 1'b1, 0, 0) c38081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38081));
	wire w39081;

	wire w42081;

	wire w43081;

	wire w46081;
	repeater #(1, 1'b1, 0, 0) c46081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46081));
	wire w47081;

	wire w40083;
	torch #(1'b0) c40083 (.i_clk(tick), .i_in(), .o_out(w40083));
	wire w26085;
	repeater #(1, 1'b0, 0, 0) c26085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26085));
	wire w27085;

	wire w30085;
	repeater #(1, 1'b0, 0, 0) c30085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30085));
	wire w31085;

	wire w34085;
	repeater #(1, 1'b1, 0, 0) c34085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34085));
	wire w35085;

	wire w38085;
	repeater #(1, 1'b0, 0, 0) c38085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38085));
	wire w39085;

	wire w42085;
	repeater #(1, 1'b1, 0, 0) c42085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42085));
	wire w43085;

	wire w46085;
	repeater #(1, 1'b0, 0, 0) c46085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46085));
	wire w47085;

	wire w50085;
	repeater #(1, 1'b0, 0, 0) c50085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50085));
	wire w51085;

	wire w26088;
	repeater #(1, 1'b0, 0, 0) c26088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26088));
	wire w31088;
	repeater #(1, 1'b0, 0, 0) c31088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31088));
	wire w34088;
	repeater #(1, 1'b1, 0, 0) c34088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34088));
	wire w39088;
	repeater #(1, 1'b0, 0, 0) c39088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39088));
	wire w42088;
	repeater #(1, 1'b1, 0, 0) c42088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42088));
	wire w47088;
	repeater #(1, 1'b0, 0, 0) c47088 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47088));
	wire w28089;

	wire w29089;

	wire w36089;

	wire w37089;

	wire w44089;

	wire w45089;

	wire w50089;
	repeater #(4, 1'b0, 0, 0) c50089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50089));
	wire w26090;
	repeater #(4, 1'b0, 0, 0) c26090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26090));
	wire w31090;
	repeater #(2, 1'b0, 0, 0) c31090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31090));
	wire w34090;
	repeater #(4, 1'b1, 0, 0) c34090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34090));
	wire w39090;
	repeater #(2, 1'b0, 0, 0) c39090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39090));
	wire w42090;
	repeater #(4, 1'b1, 0, 0) c42090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42090));
	wire w47090;
	repeater #(2, 1'b0, 0, 0) c47090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47090));
	wire w31092;
	repeater #(2, 1'b0, 0, 0) c31092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31092));
	wire w39092;
	repeater #(2, 1'b0, 0, 0) c39092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39092));
	wire w47092;
	repeater #(2, 1'b0, 0, 0) c47092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47092));
	wire w50093;
	repeater #(2, 1'b0, 0, 0) c50093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w50093));
	wire w26095;

	wire w27095;

	wire w30095;
	repeater #(1, 1'b1, 0, 0) c30095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30095));
	wire w31095;

	wire w34095;

	wire w35095;

	wire w38095;
	repeater #(1, 1'b0, 0, 0) c38095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38095));
	wire w39095;

	wire w42095;

	wire w43095;

	wire w46095;
	repeater #(1, 1'b1, 0, 0) c46095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w46095));
	wire w47095;

	wire w26098;
	repeater #(1, 1'b0, 0, 0) c26098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26098));
	wire w31098;
	repeater #(1, 1'b0, 0, 0) c31098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31098));
	wire w42098;
	repeater #(1, 1'b1, 0, 0) c42098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w42098));
	wire w47098;
	repeater #(1, 1'b0, 0, 0) c47098 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w47098));
	wire w28099;

	wire w29099;

	wire w33099;
	repeater #(1, 1'b0, 0, 0) c33099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w33099));
	wire w36099;

	wire w37099;

	wire w44099;

	wire w45099;

	wire w260100;
	repeater #(4, 1'b0, 0, 0) c260100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260100));
	wire w310100;
	repeater #(2, 1'b0, 0, 0) c310100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310100));
	wire w320100;
	repeater #(1, 1'b0, 0, 0) c320100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320100));
	wire w340100;
	repeater #(4, 1'b0, 0, 0) c340100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340100));
	wire w390100;
	repeater #(1, 1'b1, 0, 0) c390100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390100));
	wire w420100;
	repeater #(4, 1'b1, 0, 0) c420100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420100));
	wire w470100;
	repeater #(2, 1'b0, 0, 0) c470100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470100));
	wire w310102;
	repeater #(2, 1'b0, 0, 0) c310102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310102));
	wire w470102;
	repeater #(2, 1'b0, 0, 0) c470102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470102));
	wire w390103;
	repeater #(1, 1'b1, 0, 0) c390103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390103));
	wire w400103;
	repeater #(1, 1'b1, 0, 0) c400103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400103));
	wire w390104;
	repeater #(4, 1'b1, 0, 0) c390104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390104));
	wire w260105;

	wire w270105;

	wire w300105;
	repeater #(1, 1'b0, 0, 0) c300105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300105));
	wire w310105;

	wire w340105;

	wire w350105;

	wire w380105;
	repeater #(1, 1'b1, 0, 0) c380105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380105));
	wire w390105;

	wire w420105;

	wire w430105;

	wire w460105;
	repeater #(1, 1'b1, 0, 0) c460105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460105));
	wire w470105;

	wire w400107;
	torch #(1'b0) c400107 (.i_clk(tick), .i_in(), .o_out(w400107));
	wire w260109;
	repeater #(1, 1'b1, 0, 0) c260109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260109));
	wire w270109;

	wire w300109;
	repeater #(1, 1'b1, 0, 0) c300109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300109));
	wire w310109;

	wire w340109;
	repeater #(1, 1'b1, 0, 0) c340109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340109));
	wire w350109;

	wire w380109;
	repeater #(1, 1'b1, 0, 0) c380109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380109));
	wire w390109;

	wire w420109;
	repeater #(1, 1'b1, 0, 0) c420109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420109));
	wire w430109;

	wire w460109;
	repeater #(1, 1'b1, 0, 0) c460109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460109));
	wire w470109;

	wire w500109;
	repeater #(1, 1'b1, 0, 0) c500109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500109));
	wire w510109;

	wire w260112;
	repeater #(1, 1'b1, 0, 0) c260112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260112));
	wire w310112;
	repeater #(1, 1'b1, 0, 0) c310112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310112));
	wire w340112;
	repeater #(1, 1'b1, 0, 0) c340112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340112));
	wire w390112;
	repeater #(1, 1'b1, 0, 0) c390112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390112));
	wire w420112;
	repeater #(1, 1'b1, 0, 0) c420112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420112));
	wire w470112;
	repeater #(1, 1'b1, 0, 0) c470112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470112));
	wire w280113;

	wire w290113;

	wire w360113;

	wire w370113;

	wire w440113;

	wire w450113;

	wire w500113;
	repeater #(4, 1'b1, 0, 0) c500113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500113));
	wire w260114;
	repeater #(4, 1'b1, 0, 0) c260114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260114));
	wire w310114;
	repeater #(2, 1'b1, 0, 0) c310114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310114));
	wire w340114;
	repeater #(4, 1'b1, 0, 0) c340114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340114));
	wire w390114;
	repeater #(2, 1'b1, 0, 0) c390114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390114));
	wire w420114;
	repeater #(4, 1'b1, 0, 0) c420114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420114));
	wire w470114;
	repeater #(2, 1'b1, 0, 0) c470114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470114));
	wire w310116;
	repeater #(2, 1'b1, 0, 0) c310116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310116));
	wire w390116;
	repeater #(2, 1'b1, 0, 0) c390116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390116));
	wire w470116;
	repeater #(2, 1'b1, 0, 0) c470116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470116));
	wire w500117;
	repeater #(2, 1'b1, 0, 0) c500117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500117));
	wire w260119;

	wire w270119;

	wire w300119;
	repeater #(1, 1'b0, 0, 0) c300119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300119));
	wire w310119;

	wire w340119;

	wire w350119;

	wire w380119;
	repeater #(1, 1'b0, 0, 0) c380119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380119));
	wire w390119;

	wire w420119;

	wire w430119;

	wire w460119;
	repeater #(1, 1'b1, 0, 0) c460119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460119));
	wire w470119;

	wire w260122;
	repeater #(1, 1'b1, 0, 0) c260122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260122));
	wire w310122;
	repeater #(1, 1'b1, 0, 0) c310122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310122));
	wire w420122;
	repeater #(1, 1'b1, 0, 0) c420122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420122));
	wire w470122;
	repeater #(1, 1'b1, 0, 0) c470122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470122));
	wire w280123;

	wire w290123;

	wire w330123;
	repeater #(1, 1'b1, 0, 0) c330123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330123));
	wire w360123;

	wire w370123;

	wire w440123;

	wire w450123;

	wire w260124;
	repeater #(4, 1'b1, 0, 0) c260124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260124));
	wire w310124;
	repeater #(2, 1'b1, 0, 0) c310124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310124));
	wire w320124;
	repeater #(1, 1'b1, 0, 0) c320124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320124));
	wire w340124;
	repeater #(4, 1'b1, 0, 0) c340124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340124));
	wire w390124;
	repeater #(1, 1'b1, 0, 0) c390124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390124));
	wire w420124;
	repeater #(4, 1'b1, 0, 0) c420124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420124));
	wire w470124;
	repeater #(2, 1'b1, 0, 0) c470124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470124));
	wire w310126;
	repeater #(2, 1'b1, 0, 0) c310126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310126));
	wire w470126;
	repeater #(2, 1'b1, 0, 0) c470126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470126));
	wire w390127;
	repeater #(1, 1'b1, 0, 0) c390127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390127));
	wire w400127;
	repeater #(1, 1'b1, 0, 0) c400127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400127));
	wire w390128;
	repeater #(4, 1'b1, 0, 0) c390128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390128));
	wire w260129;

	wire w270129;

	wire w300129;
	repeater #(1, 1'b0, 0, 0) c300129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300129));
	wire w310129;

	wire w340129;

	wire w350129;

	wire w380129;
	repeater #(1, 1'b1, 0, 0) c380129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380129));
	wire w390129;

	wire w420129;

	wire w430129;

	wire w460129;
	repeater #(1, 1'b1, 0, 0) c460129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460129));
	wire w470129;

	wire w400131;
	torch #(1'b1) c400131 (.i_clk(tick), .i_in(), .o_out(w400131));
	wire w260133;
	repeater #(1, 1'b0, 0, 0) c260133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260133));
	wire w270133;

	wire w300133;
	repeater #(1, 1'b0, 0, 0) c300133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300133));
	wire w310133;

	wire w340133;
	repeater #(1, 1'b0, 0, 0) c340133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340133));
	wire w350133;

	wire w380133;
	repeater #(1, 1'b0, 0, 0) c380133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380133));
	wire w390133;

	wire w420133;
	repeater #(1, 1'b0, 0, 0) c420133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420133));
	wire w430133;

	wire w460133;
	repeater #(1, 1'b0, 0, 0) c460133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460133));
	wire w470133;

	wire w500133;
	repeater #(1, 1'b0, 0, 0) c500133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500133));
	wire w510133;

	wire w260136;
	repeater #(1, 1'b0, 0, 0) c260136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260136));
	wire w310136;
	repeater #(1, 1'b0, 0, 0) c310136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310136));
	wire w340136;
	repeater #(1, 1'b0, 0, 0) c340136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340136));
	wire w390136;
	repeater #(1, 1'b0, 0, 0) c390136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390136));
	wire w420136;
	repeater #(1, 1'b0, 0, 0) c420136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420136));
	wire w470136;
	repeater #(1, 1'b0, 0, 0) c470136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470136));
	wire w280137;

	wire w290137;

	wire w360137;

	wire w370137;

	wire w440137;

	wire w450137;

	wire w500137;
	repeater #(4, 1'b0, 0, 0) c500137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500137));
	wire w260138;
	repeater #(4, 1'b0, 0, 0) c260138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260138));
	wire w310138;
	repeater #(2, 1'b0, 0, 0) c310138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310138));
	wire w340138;
	repeater #(4, 1'b0, 0, 0) c340138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340138));
	wire w390138;
	repeater #(2, 1'b0, 0, 0) c390138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390138));
	wire w420138;
	repeater #(4, 1'b0, 0, 0) c420138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420138));
	wire w470138;
	repeater #(2, 1'b0, 0, 0) c470138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470138));
	wire w310140;
	repeater #(2, 1'b0, 0, 0) c310140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310140));
	wire w390140;
	repeater #(2, 1'b0, 0, 0) c390140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390140));
	wire w470140;
	repeater #(2, 1'b0, 0, 0) c470140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470140));
	wire w500141;
	repeater #(2, 1'b0, 0, 0) c500141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500141));
	wire w260143;

	wire w270143;

	wire w300143;
	repeater #(1, 1'b0, 0, 0) c300143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300143));
	wire w310143;

	wire w340143;

	wire w350143;

	wire w380143;
	repeater #(1, 1'b0, 0, 0) c380143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380143));
	wire w390143;

	wire w420143;

	wire w430143;

	wire w460143;
	repeater #(1, 1'b0, 0, 0) c460143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460143));
	wire w470143;

	wire w260146;
	repeater #(1, 1'b0, 0, 0) c260146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260146));
	wire w310146;
	repeater #(1, 1'b0, 0, 0) c310146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310146));
	wire w420146;
	repeater #(1, 1'b0, 0, 0) c420146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420146));
	wire w470146;
	repeater #(1, 1'b0, 0, 0) c470146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470146));
	wire w280147;

	wire w290147;

	wire w330147;
	repeater #(1, 1'b0, 0, 0) c330147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330147));
	wire w360147;

	wire w370147;

	wire w440147;

	wire w450147;

	wire w260148;
	repeater #(4, 1'b0, 0, 0) c260148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260148));
	wire w310148;
	repeater #(2, 1'b0, 0, 0) c310148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310148));
	wire w320148;
	repeater #(1, 1'b0, 0, 0) c320148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320148));
	wire w340148;
	repeater #(4, 1'b0, 0, 0) c340148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340148));
	wire w390148;
	repeater #(1, 1'b0, 0, 0) c390148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390148));
	wire w420148;
	repeater #(4, 1'b0, 0, 0) c420148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420148));
	wire w470148;
	repeater #(2, 1'b0, 0, 0) c470148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470148));
	wire w310150;
	repeater #(2, 1'b0, 0, 0) c310150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310150));
	wire w470150;
	repeater #(2, 1'b0, 0, 0) c470150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470150));
	wire w390151;
	repeater #(1, 1'b0, 0, 0) c390151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390151));
	wire w400151;
	repeater #(1, 1'b0, 0, 0) c400151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400151));
	wire w390152;
	repeater #(4, 1'b0, 0, 0) c390152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390152));
	wire w260153;

	wire w270153;

	wire w300153;
	repeater #(1, 1'b0, 0, 0) c300153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300153));
	wire w310153;

	wire w340153;

	wire w350153;

	wire w380153;
	repeater #(1, 1'b0, 0, 0) c380153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380153));
	wire w390153;

	wire w420153;

	wire w430153;

	wire w460153;
	repeater #(1, 1'b0, 0, 0) c460153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460153));
	wire w470153;

	wire w400155;
	torch #(1'b0) c400155 (.i_clk(tick), .i_in(), .o_out(w400155));
	wire w260157;
	repeater #(1, 1'b1, 0, 0) c260157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260157));
	wire w270157;

	wire w300157;
	repeater #(1, 1'b1, 0, 0) c300157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300157));
	wire w310157;

	wire w340157;
	repeater #(1, 1'b1, 0, 0) c340157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340157));
	wire w350157;

	wire w380157;
	repeater #(1, 1'b1, 0, 0) c380157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380157));
	wire w390157;

	wire w420157;
	repeater #(1, 1'b1, 0, 0) c420157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420157));
	wire w430157;

	wire w460157;
	repeater #(1, 1'b1, 0, 0) c460157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460157));
	wire w470157;

	wire w500157;
	repeater #(1, 1'b0, 0, 0) c500157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500157));
	wire w510157;

	wire w260160;
	repeater #(1, 1'b1, 0, 0) c260160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260160));
	wire w310160;
	repeater #(1, 1'b1, 0, 0) c310160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310160));
	wire w340160;
	repeater #(1, 1'b1, 0, 0) c340160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340160));
	wire w390160;
	repeater #(1, 1'b1, 0, 0) c390160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390160));
	wire w420160;
	repeater #(1, 1'b1, 0, 0) c420160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420160));
	wire w470160;
	repeater #(1, 1'b1, 0, 0) c470160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470160));
	wire w280161;

	wire w290161;

	wire w360161;

	wire w370161;

	wire w440161;

	wire w450161;

	wire w500161;
	repeater #(4, 1'b0, 0, 0) c500161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500161));
	wire w260162;
	repeater #(4, 1'b1, 0, 0) c260162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260162));
	wire w310162;
	repeater #(2, 1'b1, 0, 0) c310162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310162));
	wire w340162;
	repeater #(4, 1'b1, 0, 0) c340162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340162));
	wire w390162;
	repeater #(2, 1'b1, 0, 0) c390162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390162));
	wire w420162;
	repeater #(4, 1'b1, 0, 0) c420162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420162));
	wire w470162;
	repeater #(2, 1'b1, 0, 0) c470162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470162));
	wire w310164;
	repeater #(2, 1'b1, 0, 0) c310164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310164));
	wire w390164;
	repeater #(2, 1'b1, 0, 0) c390164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390164));
	wire w470164;
	repeater #(2, 1'b1, 0, 0) c470164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470164));
	wire w500165;
	repeater #(2, 1'b0, 0, 0) c500165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w500165));
	wire w260167;

	wire w270167;

	wire w300167;
	repeater #(1, 1'b0, 0, 0) c300167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300167));
	wire w310167;

	wire w340167;

	wire w350167;

	wire w380167;
	repeater #(1, 1'b0, 0, 0) c380167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380167));
	wire w390167;

	wire w420167;

	wire w430167;

	wire w460167;
	repeater #(1, 1'b0, 0, 0) c460167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460167));
	wire w470167;

	wire w260170;
	repeater #(1, 1'b1, 0, 0) c260170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260170));
	wire w310170;
	repeater #(1, 1'b1, 0, 0) c310170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310170));
	wire w420170;
	repeater #(1, 1'b1, 0, 0) c420170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420170));
	wire w470170;
	repeater #(1, 1'b0, 0, 0) c470170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470170));
	wire w280171;

	wire w290171;

	wire w330171;
	repeater #(1, 1'b1, 0, 0) c330171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w330171));
	wire w360171;

	wire w370171;

	wire w440171;

	wire w450171;

	wire w260172;
	repeater #(4, 1'b1, 0, 0) c260172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260172));
	wire w310172;
	repeater #(2, 1'b1, 0, 0) c310172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310172));
	wire w320172;
	repeater #(1, 1'b1, 0, 0) c320172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w320172));
	wire w340172;
	repeater #(4, 1'b1, 0, 0) c340172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340172));
	wire w390172;
	repeater #(1, 1'b1, 0, 0) c390172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390172));
	wire w420172;
	repeater #(4, 1'b1, 0, 0) c420172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w420172));
	wire w470172;
	repeater #(2, 1'b0, 0, 0) c470172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470172));
	wire w310174;
	repeater #(2, 1'b1, 0, 0) c310174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310174));
	wire w470174;
	repeater #(2, 1'b0, 0, 0) c470174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w470174));
	wire w390175;
	repeater #(1, 1'b1, 0, 0) c390175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390175));
	wire w400175;
	repeater #(1, 1'b1, 0, 0) c400175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w400175));
	wire w390176;
	repeater #(4, 1'b1, 0, 0) c390176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w390176));
	wire w260177;

	wire w270177;

	wire w300177;
	repeater #(1, 1'b0, 0, 0) c300177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300177));
	wire w310177;

	wire w340177;

	wire w350177;

	wire w380177;
	repeater #(1, 1'b0, 0, 0) c380177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w380177));
	wire w390177;

	wire w420177;

	wire w430177;

	wire w460177;
	repeater #(1, 1'b1, 0, 0) c460177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w460177));
	wire w470177;

	wire w4010;
	torch #(1'b1) c4010 (.i_clk(tick), .i_in(), .o_out(w4010));
	wire w25154;
	repeater #(1, 1'b0, 0, 0) c25154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25154));
	wire w26155;
	repeater #(1, 1'b0, 0, 0) c26155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26155));
	wire w196155;
	repeater #(1, 1'b1, 0, 0) c196155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196155));
	wire w5156;
	repeater #(2, 1'b1, 0, 0) c5156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w5156));
	wire w6156;
	repeater #(1, 1'b1, 0, 0) c6156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6156));
	wire w7156;

	wire w22156;

	wire w25156;
	repeater #(1, 1'b1, 0, 0) c25156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w25156));
	wire w35156;
	repeater #(1, 1'b1, 0, 0) c35156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w35156));
	wire w40156;
	repeater #(1, 1'b1, 0, 0) c40156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40156));
	wire w24157;
	repeater #(1, 1'b0, 0, 0) c24157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24157));
	wire w37157;

	wire w38157;

	wire w38159;
	repeater #(1, 1'b0, 0, 0) c38159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38159));
	wire w52159;
	repeater #(1, 1'b1, 0, 0) c52159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52159));
	wire w52160;

	wire w54161;
	repeater #(1, 1'b0, 0, 0) c54161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54161));
	wire w23162;
	repeater #(1, 1'b0, 0, 0) c23162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23162));
	wire w193169;
	repeater #(1, 1'b0, 0, 0) c193169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193169));
	wire w54177;
	repeater #(1, 1'b0, 0, 0) c54177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54177));
	wire w52183;
	repeater #(1, 1'b1, 0, 0) c52183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w52183));
	wire w52184;

	wire w54185;
	repeater #(1, 1'b0, 0, 0) c54185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w54185));
	wire w541101;
	repeater #(1, 1'b0, 0, 0) c541101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w541101));
	wire w521107;
	repeater #(1, 1'b1, 0, 0) c521107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w521107));
	wire w521108;

	wire w541109;
	repeater #(1, 1'b0, 0, 0) c541109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w541109));
	wire w541125;
	repeater #(1, 1'b0, 0, 0) c541125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w541125));
	wire w521131;
	repeater #(1, 1'b1, 0, 0) c521131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w521131));
	wire w521132;

	wire w541133;
	repeater #(1, 1'b0, 0, 0) c541133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w541133));
	wire w38013;
	repeater #(1, 1'b0, 0, 0) c38013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38013));
	wire w36019;
	repeater #(1, 1'b1, 0, 0) c36019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w36019));
	wire w36020;

	wire w38021;
	repeater #(1, 1'b0, 0, 0) c38021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38021));
	wire w38037;
	repeater #(1, 1'b0, 0, 0) c38037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w38037));
	wire w40042;
	repeater #(1, 1'b0, 0, 0) c40042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40042));
	wire w41044;

	wire w44044;
	assign outputs[120] = ();
	wire w41045;

	wire w39046;
	repeater #(1, 1'b0, 0, 0) c39046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w39046));
	wire w181098;

	wire w100104;
	repeater #(1, 1'b0, 0, 0) c100104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100104));
	wire w110104;

	wire w140104;
	repeater #(1, 1'b1, 0, 0) c140104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140104));
	wire w150104;

	wire w180104;
	repeater #(1, 1'b1, 0, 0) c180104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180104));
	wire w190104;

	wire w220104;
	repeater #(1, 1'b0, 0, 0) c220104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220104));
	wire w230104;

	wire w260104;
	repeater #(1, 1'b0, 0, 0) c260104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260104));
	wire w270104;

	wire w300104;
	repeater #(1, 1'b1, 0, 0) c300104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300104));
	wire w310104;

	wire w340104;
	repeater #(1, 1'b1, 0, 0) c340104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340104));
	wire w350104;

	wire w100107;
	repeater #(1, 1'b0, 0, 0) c100107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100107));
	wire w150107;
	repeater #(1, 1'b1, 0, 0) c150107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150107));
	wire w180107;
	repeater #(1, 1'b1, 0, 0) c180107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180107));
	wire w230107;
	repeater #(1, 1'b0, 0, 0) c230107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230107));
	wire w260107;
	repeater #(1, 1'b0, 0, 0) c260107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260107));
	wire w310107;
	repeater #(1, 1'b1, 0, 0) c310107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310107));
	wire w120108;

	wire w130108;

	wire w200108;

	wire w210108;

	wire w280108;

	wire w290108;

	wire w340108;
	repeater #(4, 1'b1, 0, 0) c340108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340108));
	wire w100109;
	repeater #(4, 1'b0, 0, 0) c100109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100109));
	wire w150109;
	repeater #(2, 1'b1, 0, 0) c150109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150109));
	wire w180109;
	repeater #(4, 1'b1, 0, 0) c180109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180109));
	wire w230109;
	repeater #(2, 1'b0, 0, 0) c230109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230109));
	wire w260109;
	repeater #(4, 1'b0, 0, 0) c260109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260109));
	wire w310109;
	repeater #(2, 1'b1, 0, 0) c310109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310109));
	wire w150111;
	repeater #(2, 1'b1, 0, 0) c150111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150111));
	wire w230111;
	repeater #(2, 1'b0, 0, 0) c230111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230111));
	wire w310111;
	repeater #(2, 1'b1, 0, 0) c310111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310111));
	wire w1780111;

	wire w340112;
	repeater #(2, 1'b1, 0, 0) c340112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340112));
	wire w100114;

	wire w110114;

	wire w140114;
	repeater #(1, 1'b0, 0, 0) c140114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140114));
	wire w150114;

	wire w180114;

	wire w190114;

	wire w220114;
	repeater #(1, 1'b1, 0, 0) c220114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220114));
	wire w230114;

	wire w260114;

	wire w270114;

	wire w300114;
	repeater #(1, 1'b1, 0, 0) c300114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300114));
	wire w310114;

	wire w100117;
	repeater #(1, 1'b1, 0, 0) c100117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100117));
	wire w150117;
	repeater #(1, 1'b1, 0, 0) c150117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150117));
	wire w260117;
	repeater #(1, 1'b0, 0, 0) c260117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260117));
	wire w310117;
	repeater #(1, 1'b1, 0, 0) c310117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310117));
	wire w120118;

	wire w130118;

	wire w170118;
	repeater #(1, 1'b1, 0, 0) c170118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170118));
	wire w200118;

	wire w210118;

	wire w280118;

	wire w290118;

	wire w100119;
	repeater #(4, 1'b1, 0, 0) c100119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100119));
	wire w150119;
	repeater #(2, 1'b1, 0, 0) c150119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150119));
	wire w160119;
	repeater #(1, 1'b1, 0, 0) c160119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160119));
	wire w180119;
	repeater #(4, 1'b1, 0, 0) c180119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180119));
	wire w230119;
	repeater #(1, 1'b0, 0, 0) c230119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230119));
	wire w260119;
	repeater #(4, 1'b0, 0, 0) c260119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260119));
	wire w310119;
	repeater #(2, 1'b1, 0, 0) c310119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310119));
	wire w150121;
	repeater #(2, 1'b1, 0, 0) c150121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150121));
	wire w310121;
	repeater #(2, 1'b1, 0, 0) c310121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310121));
	wire w230122;
	repeater #(1, 1'b0, 0, 0) c230122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230122));
	wire w240122;
	repeater #(1, 1'b0, 0, 0) c240122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240122));
	wire w230123;
	repeater #(4, 1'b0, 0, 0) c230123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230123));
	wire w100124;

	wire w110124;

	wire w140124;
	repeater #(1, 1'b0, 0, 0) c140124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140124));
	wire w150124;

	wire w180124;

	wire w190124;

	wire w220124;
	repeater #(1, 1'b1, 0, 0) c220124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220124));
	wire w230124;

	wire w260124;

	wire w270124;

	wire w300124;
	repeater #(1, 1'b1, 0, 0) c300124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300124));
	wire w310124;

	wire w240126;
	torch #(1'b1) c240126 (.i_clk(tick), .i_in(), .o_out(w240126));
	wire w100128;
	repeater #(1, 1'b1, 0, 0) c100128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100128));
	wire w110128;

	wire w140128;
	repeater #(1, 1'b1, 0, 0) c140128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140128));
	wire w150128;

	wire w180128;
	repeater #(1, 1'b1, 0, 0) c180128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180128));
	wire w190128;

	wire w220128;
	repeater #(1, 1'b1, 0, 0) c220128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220128));
	wire w230128;

	wire w260128;
	repeater #(1, 1'b1, 0, 0) c260128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260128));
	wire w270128;

	wire w300128;
	repeater #(1, 1'b1, 0, 0) c300128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300128));
	wire w310128;

	wire w340128;
	repeater #(1, 1'b1, 0, 0) c340128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340128));
	wire w350128;

	wire w100131;
	repeater #(1, 1'b1, 0, 0) c100131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100131));
	wire w150131;
	repeater #(1, 1'b1, 0, 0) c150131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150131));
	wire w180131;
	repeater #(1, 1'b1, 0, 0) c180131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180131));
	wire w230131;
	repeater #(1, 1'b1, 0, 0) c230131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230131));
	wire w260131;
	repeater #(1, 1'b1, 0, 0) c260131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260131));
	wire w310131;
	repeater #(1, 1'b1, 0, 0) c310131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310131));
	wire w120132;

	wire w130132;

	wire w200132;

	wire w210132;

	wire w280132;

	wire w290132;

	wire w340132;
	repeater #(4, 1'b1, 0, 0) c340132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340132));
	wire w100133;
	repeater #(4, 1'b1, 0, 0) c100133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100133));
	wire w150133;
	repeater #(2, 1'b1, 0, 0) c150133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150133));
	wire w180133;
	repeater #(4, 1'b1, 0, 0) c180133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180133));
	wire w230133;
	repeater #(2, 1'b1, 0, 0) c230133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230133));
	wire w260133;
	repeater #(4, 1'b1, 0, 0) c260133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260133));
	wire w310133;
	repeater #(2, 1'b1, 0, 0) c310133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310133));
	wire w150135;
	repeater #(2, 1'b1, 0, 0) c150135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150135));
	wire w230135;
	repeater #(2, 1'b1, 0, 0) c230135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230135));
	wire w310135;
	repeater #(2, 1'b1, 0, 0) c310135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310135));
	wire w340136;
	repeater #(2, 1'b1, 0, 0) c340136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340136));
	wire w100138;

	wire w110138;

	wire w140138;
	repeater #(1, 1'b1, 0, 0) c140138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140138));
	wire w150138;

	wire w180138;

	wire w190138;

	wire w220138;
	repeater #(1, 1'b0, 0, 0) c220138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220138));
	wire w230138;

	wire w260138;

	wire w270138;

	wire w300138;
	repeater #(1, 1'b1, 0, 0) c300138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300138));
	wire w310138;

	wire w100141;
	repeater #(1, 1'b1, 0, 0) c100141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100141));
	wire w150141;
	repeater #(1, 1'b1, 0, 0) c150141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150141));
	wire w260141;
	repeater #(1, 1'b1, 0, 0) c260141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260141));
	wire w310141;
	repeater #(1, 1'b1, 0, 0) c310141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310141));
	wire w120142;

	wire w130142;

	wire w170142;
	repeater #(1, 1'b1, 0, 0) c170142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170142));
	wire w200142;

	wire w210142;

	wire w280142;

	wire w290142;

	wire w100143;
	repeater #(4, 1'b1, 0, 0) c100143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100143));
	wire w150143;
	repeater #(2, 1'b1, 0, 0) c150143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150143));
	wire w160143;
	repeater #(1, 1'b1, 0, 0) c160143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160143));
	wire w180143;
	repeater #(4, 1'b1, 0, 0) c180143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180143));
	wire w230143;
	repeater #(1, 1'b1, 0, 0) c230143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230143));
	wire w260143;
	repeater #(4, 1'b1, 0, 0) c260143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260143));
	wire w310143;
	repeater #(2, 1'b1, 0, 0) c310143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310143));
	wire w150145;
	repeater #(2, 1'b1, 0, 0) c150145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150145));
	wire w310145;
	repeater #(2, 1'b1, 0, 0) c310145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310145));
	wire w230146;
	repeater #(1, 1'b1, 0, 0) c230146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230146));
	wire w240146;
	repeater #(1, 1'b1, 0, 0) c240146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240146));
	wire w230147;
	repeater #(4, 1'b1, 0, 0) c230147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230147));
	wire w100148;

	wire w110148;

	wire w140148;
	repeater #(1, 1'b0, 0, 0) c140148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140148));
	wire w150148;

	wire w180148;

	wire w190148;

	wire w220148;
	repeater #(1, 1'b1, 0, 0) c220148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220148));
	wire w230148;

	wire w260148;

	wire w270148;

	wire w300148;
	repeater #(1, 1'b1, 0, 0) c300148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300148));
	wire w310148;

	wire w240150;
	torch #(1'b1) c240150 (.i_clk(tick), .i_in(), .o_out(w240150));
	wire w100152;
	repeater #(1, 1'b0, 0, 0) c100152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100152));
	wire w110152;

	wire w140152;
	repeater #(1, 1'b0, 0, 0) c140152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140152));
	wire w150152;

	wire w180152;
	repeater #(1, 1'b1, 0, 0) c180152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180152));
	wire w190152;

	wire w220152;
	repeater #(1, 1'b0, 0, 0) c220152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220152));
	wire w230152;

	wire w260152;
	repeater #(1, 1'b1, 0, 0) c260152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260152));
	wire w270152;

	wire w300152;
	repeater #(1, 1'b0, 0, 0) c300152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300152));
	wire w310152;

	wire w340152;
	repeater #(1, 1'b0, 0, 0) c340152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340152));
	wire w350152;

	wire w100155;
	repeater #(1, 1'b0, 0, 0) c100155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100155));
	wire w150155;
	repeater #(1, 1'b0, 0, 0) c150155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150155));
	wire w180155;
	repeater #(1, 1'b1, 0, 0) c180155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180155));
	wire w230155;
	repeater #(1, 1'b0, 0, 0) c230155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230155));
	wire w260155;
	repeater #(1, 1'b1, 0, 0) c260155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260155));
	wire w310155;
	repeater #(1, 1'b0, 0, 0) c310155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310155));
	wire w120156;

	wire w130156;

	wire w200156;

	wire w210156;

	wire w280156;

	wire w290156;

	wire w340156;
	repeater #(4, 1'b0, 0, 0) c340156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340156));
	wire w100157;
	repeater #(4, 1'b0, 0, 0) c100157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100157));
	wire w150157;
	repeater #(2, 1'b0, 0, 0) c150157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150157));
	wire w180157;
	repeater #(4, 1'b1, 0, 0) c180157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180157));
	wire w230157;
	repeater #(2, 1'b0, 0, 0) c230157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230157));
	wire w260157;
	repeater #(4, 1'b1, 0, 0) c260157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260157));
	wire w310157;
	repeater #(2, 1'b0, 0, 0) c310157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310157));
	wire w150159;
	repeater #(2, 1'b0, 0, 0) c150159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150159));
	wire w230159;
	repeater #(2, 1'b0, 0, 0) c230159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230159));
	wire w310159;
	repeater #(2, 1'b0, 0, 0) c310159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310159));
	wire w340160;
	repeater #(2, 1'b0, 0, 0) c340160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340160));
	wire w100162;

	wire w110162;

	wire w140162;
	repeater #(1, 1'b0, 0, 0) c140162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140162));
	wire w150162;

	wire w180162;

	wire w190162;

	wire w220162;
	repeater #(1, 1'b0, 0, 0) c220162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220162));
	wire w230162;

	wire w260162;

	wire w270162;

	wire w300162;
	repeater #(1, 1'b1, 0, 0) c300162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300162));
	wire w310162;

	wire w100165;
	repeater #(1, 1'b0, 0, 0) c100165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100165));
	wire w150165;
	repeater #(1, 1'b0, 0, 0) c150165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150165));
	wire w260165;
	repeater #(1, 1'b1, 0, 0) c260165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260165));
	wire w310165;
	repeater #(1, 1'b0, 0, 0) c310165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310165));
	wire w120166;

	wire w130166;

	wire w170166;
	repeater #(1, 1'b0, 0, 0) c170166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170166));
	wire w200166;

	wire w210166;

	wire w280166;

	wire w290166;

	wire w100167;
	repeater #(4, 1'b0, 0, 0) c100167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100167));
	wire w150167;
	repeater #(2, 1'b0, 0, 0) c150167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150167));
	wire w160167;
	repeater #(1, 1'b0, 0, 0) c160167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160167));
	wire w180167;
	repeater #(4, 1'b0, 0, 0) c180167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180167));
	wire w230167;
	repeater #(1, 1'b1, 0, 0) c230167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230167));
	wire w260167;
	repeater #(4, 1'b1, 0, 0) c260167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260167));
	wire w310167;
	repeater #(2, 1'b0, 0, 0) c310167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310167));
	wire w150169;
	repeater #(2, 1'b0, 0, 0) c150169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150169));
	wire w310169;
	repeater #(2, 1'b0, 0, 0) c310169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w310169));
	wire w230170;
	repeater #(1, 1'b1, 0, 0) c230170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230170));
	wire w240170;
	repeater #(1, 1'b1, 0, 0) c240170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w240170));
	wire w230171;
	repeater #(4, 1'b1, 0, 0) c230171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w230171));
	wire w100172;

	wire w110172;

	wire w140172;
	repeater #(1, 1'b0, 0, 0) c140172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140172));
	wire w150172;

	wire w180172;

	wire w190172;

	wire w220172;
	repeater #(1, 1'b1, 0, 0) c220172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220172));
	wire w230172;

	wire w260172;

	wire w270172;

	wire w300172;
	repeater #(1, 1'b1, 0, 0) c300172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300172));
	wire w310172;

	wire w240174;
	torch #(1'b0) c240174 (.i_clk(tick), .i_in(), .o_out(w240174));
	wire w100176;
	repeater #(1, 1'b0, 0, 0) c100176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100176));
	wire w110176;

	wire w140176;
	repeater #(1, 1'b0, 0, 0) c140176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140176));
	wire w150176;

	wire w180176;
	repeater #(1, 1'b0, 0, 0) c180176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180176));
	wire w190176;

	wire w220176;
	repeater #(1, 1'b0, 0, 0) c220176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w220176));
	wire w230176;

	wire w260176;
	repeater #(1, 1'b0, 0, 0) c260176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w260176));
	wire w270176;

	wire w300176;
	repeater #(1, 1'b0, 0, 0) c300176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w300176));
	wire w310176;

	wire w340176;
	repeater #(1, 1'b0, 0, 0) c340176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w340176));
	wire w350176;

	wire w1010;
	repeater #(1, 1'b0, 0, 0) c1010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1010));
	wire w1510;
	repeater #(1, 1'b0, 0, 0) c1510 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1510));
	wire w1810;
	repeater #(1, 1'b0, 0, 0) c1810 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810));
	wire w2310;
	repeater #(1, 1'b0, 0, 0) c2310 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2310));
	wire w2610;
	repeater #(1, 1'b0, 0, 0) c2610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2610));
	wire w3110;
	repeater #(1, 1'b0, 0, 0) c3110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3110));
	wire w1211;

	wire w1311;

	wire w2011;

	wire w2111;

	wire w2811;

	wire w2911;

	wire w3411;
	repeater #(4, 1'b0, 0, 0) c3411 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3411));
	wire w1012;
	repeater #(4, 1'b0, 0, 0) c1012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1012));
	wire w1512;
	repeater #(2, 1'b0, 0, 0) c1512 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1512));
	wire w1812;
	repeater #(4, 1'b0, 0, 0) c1812 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1812));
	wire w2312;
	repeater #(2, 1'b0, 0, 0) c2312 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2312));
	wire w2612;
	repeater #(4, 1'b0, 0, 0) c2612 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2612));
	wire w3112;
	repeater #(2, 1'b0, 0, 0) c3112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3112));
	wire w1514;
	repeater #(2, 1'b0, 0, 0) c1514 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1514));
	wire w2314;
	repeater #(2, 1'b0, 0, 0) c2314 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2314));
	wire w3114;
	repeater #(2, 1'b0, 0, 0) c3114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3114));
	wire w3415;
	repeater #(2, 1'b0, 0, 0) c3415 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3415));
	wire w1017;

	wire w1117;

	wire w1417;
	repeater #(1, 1'b0, 0, 0) c1417 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1417));
	wire w1517;

	wire w1817;

	wire w1917;

	wire w2217;
	repeater #(1, 1'b0, 0, 0) c2217 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2217));
	wire w2317;

	wire w2617;

	wire w2717;

	wire w3017;
	repeater #(1, 1'b0, 0, 0) c3017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w3017));
	wire w3117;

	wire w10110;
	repeater #(1, 1'b0, 0, 0) c10110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10110));
	wire w15110;
	repeater #(1, 1'b0, 0, 0) c15110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15110));
	wire w26110;
	repeater #(1, 1'b0, 0, 0) c26110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26110));
	wire w31110;
	repeater #(1, 1'b0, 0, 0) c31110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31110));
	wire w12111;

	wire w13111;

	wire w17111;
	repeater #(1, 1'b0, 0, 0) c17111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17111));
	wire w20111;

	wire w21111;

	wire w28111;

	wire w29111;

	wire w10112;
	repeater #(4, 1'b0, 0, 0) c10112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10112));
	wire w15112;
	repeater #(2, 1'b0, 0, 0) c15112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15112));
	wire w16112;
	repeater #(1, 1'b0, 0, 0) c16112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16112));
	wire w18112;
	repeater #(4, 1'b0, 0, 0) c18112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18112));
	wire w23112;
	repeater #(1, 1'b0, 0, 0) c23112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23112));
	wire w26112;
	repeater #(4, 1'b0, 0, 0) c26112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26112));
	wire w31112;
	repeater #(2, 1'b0, 0, 0) c31112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31112));
	wire w15114;
	repeater #(2, 1'b0, 0, 0) c15114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15114));
	wire w31114;
	repeater #(2, 1'b0, 0, 0) c31114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31114));
	wire w23115;
	repeater #(1, 1'b0, 0, 0) c23115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23115));
	wire w24115;
	repeater #(1, 1'b0, 0, 0) c24115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24115));
	wire w23116;
	repeater #(4, 1'b0, 0, 0) c23116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23116));
	wire w10117;

	wire w11117;

	wire w14117;
	repeater #(1, 1'b0, 0, 0) c14117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14117));
	wire w15117;

	wire w18117;

	wire w19117;

	wire w22117;
	repeater #(1, 1'b0, 0, 0) c22117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22117));
	wire w23117;

	wire w26117;

	wire w27117;

	wire w30117;
	repeater #(1, 1'b0, 0, 0) c30117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30117));
	wire w31117;

	wire w24119;
	torch #(1'b0) c24119 (.i_clk(tick), .i_in(), .o_out(w24119));
	wire w10121;
	repeater #(1, 1'b1, 0, 0) c10121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10121));
	wire w11121;

	wire w14121;
	repeater #(1, 1'b1, 0, 0) c14121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14121));
	wire w15121;

	wire w18121;
	repeater #(1, 1'b1, 0, 0) c18121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18121));
	wire w19121;

	wire w22121;
	repeater #(1, 1'b1, 0, 0) c22121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22121));
	wire w23121;

	wire w26121;
	repeater #(1, 1'b1, 0, 0) c26121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26121));
	wire w27121;

	wire w30121;
	repeater #(1, 1'b1, 0, 0) c30121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30121));
	wire w31121;

	wire w34121;
	repeater #(1, 1'b0, 0, 0) c34121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34121));
	wire w35121;

	wire w10124;
	repeater #(1, 1'b1, 0, 0) c10124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10124));
	wire w15124;
	repeater #(1, 1'b1, 0, 0) c15124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15124));
	wire w18124;
	repeater #(1, 1'b1, 0, 0) c18124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18124));
	wire w23124;
	repeater #(1, 1'b1, 0, 0) c23124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23124));
	wire w26124;
	repeater #(1, 1'b1, 0, 0) c26124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26124));
	wire w31124;
	repeater #(1, 1'b1, 0, 0) c31124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31124));
	wire w12125;

	wire w13125;

	wire w20125;

	wire w21125;

	wire w28125;

	wire w29125;

	wire w34125;
	repeater #(4, 1'b0, 0, 0) c34125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34125));
	wire w10126;
	repeater #(4, 1'b1, 0, 0) c10126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10126));
	wire w15126;
	repeater #(2, 1'b1, 0, 0) c15126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15126));
	wire w18126;
	repeater #(4, 1'b1, 0, 0) c18126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18126));
	wire w23126;
	repeater #(2, 1'b1, 0, 0) c23126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23126));
	wire w26126;
	repeater #(4, 1'b1, 0, 0) c26126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26126));
	wire w31126;
	repeater #(2, 1'b1, 0, 0) c31126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31126));
	wire w15128;
	repeater #(2, 1'b1, 0, 0) c15128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15128));
	wire w23128;
	repeater #(2, 1'b1, 0, 0) c23128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23128));
	wire w31128;
	repeater #(2, 1'b1, 0, 0) c31128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31128));
	wire w34129;
	repeater #(2, 1'b0, 0, 0) c34129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w34129));
	wire w10131;

	wire w11131;

	wire w14131;
	repeater #(1, 1'b0, 0, 0) c14131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14131));
	wire w15131;

	wire w18131;

	wire w19131;

	wire w22131;
	repeater #(1, 1'b0, 0, 0) c22131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22131));
	wire w23131;

	wire w26131;

	wire w27131;

	wire w30131;
	repeater #(1, 1'b0, 0, 0) c30131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30131));
	wire w31131;

	wire w10134;
	repeater #(1, 1'b1, 0, 0) c10134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10134));
	wire w15134;
	repeater #(1, 1'b1, 0, 0) c15134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15134));
	wire w26134;
	repeater #(1, 1'b1, 0, 0) c26134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26134));
	wire w31134;
	repeater #(1, 1'b0, 0, 0) c31134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31134));
	wire w12135;

	wire w13135;

	wire w17135;
	repeater #(1, 1'b1, 0, 0) c17135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17135));
	wire w20135;

	wire w21135;

	wire w28135;

	wire w29135;

	wire w10136;
	repeater #(4, 1'b1, 0, 0) c10136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10136));
	wire w15136;
	repeater #(2, 1'b1, 0, 0) c15136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15136));
	wire w16136;
	repeater #(1, 1'b1, 0, 0) c16136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16136));
	wire w18136;
	repeater #(4, 1'b1, 0, 0) c18136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18136));
	wire w23136;
	repeater #(1, 1'b1, 0, 0) c23136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23136));
	wire w26136;
	repeater #(4, 1'b1, 0, 0) c26136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w26136));
	wire w31136;
	repeater #(2, 1'b0, 0, 0) c31136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31136));
	wire w15138;
	repeater #(2, 1'b1, 0, 0) c15138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15138));
	wire w31138;
	repeater #(2, 1'b0, 0, 0) c31138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w31138));
	wire w23139;
	repeater #(1, 1'b1, 0, 0) c23139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23139));
	wire w24139;
	repeater #(1, 1'b1, 0, 0) c24139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24139));
	wire w23140;
	repeater #(4, 1'b1, 0, 0) c23140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23140));
	wire w10141;

	wire w11141;

	wire w14141;
	repeater #(1, 1'b0, 0, 0) c14141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14141));
	wire w15141;

	wire w18141;

	wire w19141;

	wire w22141;
	repeater #(1, 1'b0, 0, 0) c22141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22141));
	wire w23141;

	wire w26141;

	wire w27141;

	wire w30141;
	repeater #(1, 1'b1, 0, 0) c30141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w30141));
	wire w31141;

	wire w24143;
	torch #(1'b1) c24143 (.i_clk(tick), .i_in(), .o_out(w24143));
	wire w9197;
	repeater #(1, 1'b0, 0, 0) c9197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9197));
	wire w10198;
	repeater #(1, 1'b0, 0, 0) c10198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10198));
	wire w180198;
	repeater #(1, 1'b0, 0, 0) c180198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180198));
	wire w197198;
	repeater #(2, 1'b0, 0, 0) c197198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w197198));
	wire w198198;
	repeater #(1, 1'b0, 0, 0) c198198 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198198));
	wire w199198;

	wire w6199;

	wire w9199;
	repeater #(1, 1'b0, 0, 0) c9199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9199));
	wire w19199;
	repeater #(1, 1'b0, 0, 0) c19199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19199));
	wire w24199;
	repeater #(1, 1'b1, 0, 0) c24199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24199));
	wire w81100;
	repeater #(1, 1'b0, 0, 0) c81100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w81100));
	wire w211100;

	wire w221100;

	wire w221102;
	repeater #(1, 1'b1, 0, 0) c221102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w221102));
	wire w361102;
	repeater #(1, 1'b1, 0, 0) c361102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w361102));
	wire w361103;

	wire w381104;
	repeater #(1, 1'b0, 0, 0) c381104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w381104));
	wire w71105;
	repeater #(1, 1'b0, 0, 0) c71105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w71105));
	wire w1781112;
	repeater #(1, 1'b1, 0, 0) c1781112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781112));
	wire w381120;
	repeater #(1, 1'b0, 0, 0) c381120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w381120));
	wire w361126;
	repeater #(1, 1'b1, 0, 0) c361126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w361126));
	wire w361127;

	wire w381128;
	repeater #(1, 1'b0, 0, 0) c381128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w381128));
	wire w2208;
	repeater #(1, 1'b0, 0, 0) c2208 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2208));
	wire w20014;
	repeater #(1, 1'b1, 0, 0) c20014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20014));
	wire w20015;

	wire w22016;
	repeater #(1, 1'b0, 0, 0) c22016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22016));
	wire w22032;
	repeater #(1, 1'b0, 0, 0) c22032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22032));
	wire w20038;
	repeater #(1, 1'b1, 0, 0) c20038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20038));
	wire w20039;

	wire w22040;
	repeater #(1, 1'b0, 0, 0) c22040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22040));
	wire w22056;
	repeater #(1, 1'b0, 0, 0) c22056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22056));
	wire w20062;
	repeater #(1, 1'b1, 0, 0) c20062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20062));
	wire w20063;

	wire w22064;
	repeater #(1, 1'b0, 0, 0) c22064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22064));
	wire w22080;
	repeater #(1, 1'b0, 0, 0) c22080 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w22080));
	wire w24085;
	repeater #(1, 1'b0, 0, 0) c24085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w24085));
	wire w25087;

	wire w28087;
	assign outputs[121] = ();
	wire w25088;

	wire w23089;
	repeater #(1, 1'b0, 0, 0) c23089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w23089));
	wire w1650141;

	wire w2020146;
	repeater #(1, 1'b1, 0, 0) c2020146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020146));
	wire w2030146;

	wire w2060146;
	repeater #(1, 1'b1, 0, 0) c2060146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060146));
	wire w2070146;

	wire w20147;
	repeater #(1, 1'b1, 0, 0) c20147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20147));
	wire w30147;

	wire w60147;
	repeater #(1, 1'b1, 0, 0) c60147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60147));
	wire w70147;

	wire w100147;
	repeater #(1, 1'b0, 0, 0) c100147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100147));
	wire w110147;

	wire w140147;
	repeater #(1, 1'b1, 0, 0) c140147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140147));
	wire w150147;

	wire w180147;
	repeater #(1, 1'b1, 0, 0) c180147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180147));
	wire w190147;

	wire w2020149;
	repeater #(1, 1'b1, 0, 0) c2020149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020149));
	wire w2070149;
	repeater #(1, 1'b1, 0, 0) c2070149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070149));
	wire w20150;
	repeater #(1, 1'b1, 0, 0) c20150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20150));
	wire w70150;
	repeater #(1, 1'b1, 0, 0) c70150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70150));
	wire w100150;
	repeater #(1, 1'b0, 0, 0) c100150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100150));
	wire w150150;
	repeater #(1, 1'b1, 0, 0) c150150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150150));
	wire w2040150;

	wire w2050150;

	wire w40151;

	wire w50151;

	wire w120151;

	wire w130151;

	wire w180151;
	repeater #(4, 1'b1, 0, 0) c180151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180151));
	wire w2020151;
	repeater #(4, 1'b1, 0, 0) c2020151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020151));
	wire w2070151;
	repeater #(2, 1'b1, 0, 0) c2070151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070151));
	wire w20152;
	repeater #(4, 1'b1, 0, 0) c20152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20152));
	wire w70152;
	repeater #(2, 1'b1, 0, 0) c70152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70152));
	wire w100152;
	repeater #(4, 1'b0, 0, 0) c100152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100152));
	wire w150152;
	repeater #(2, 1'b1, 0, 0) c150152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150152));
	wire w2070153;
	repeater #(2, 1'b1, 0, 0) c2070153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070153));
	wire w70154;
	repeater #(2, 1'b1, 0, 0) c70154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70154));
	wire w150154;
	repeater #(2, 1'b1, 0, 0) c150154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150154));
	wire w1610154;

	wire w180155;
	repeater #(2, 1'b1, 0, 0) c180155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180155));
	wire w2020156;

	wire w2030156;

	wire w2060156;
	repeater #(1, 1'b0, 0, 0) c2060156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060156));
	wire w2070156;

	wire w20157;

	wire w30157;

	wire w60157;
	repeater #(1, 1'b1, 0, 0) c60157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60157));
	wire w70157;

	wire w100157;

	wire w110157;

	wire w140157;
	repeater #(1, 1'b1, 0, 0) c140157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140157));
	wire w150157;

	wire w2020159;
	repeater #(1, 1'b1, 0, 0) c2020159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020159));
	wire w2070159;
	repeater #(1, 1'b1, 0, 0) c2070159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070159));
	wire w100160;
	repeater #(1, 1'b0, 0, 0) c100160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100160));
	wire w150160;
	repeater #(1, 1'b1, 0, 0) c150160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150160));
	wire w2040160;

	wire w2050160;

	wire w10161;
	repeater #(1, 1'b1, 0, 0) c10161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10161));
	wire w40161;

	wire w50161;

	wire w120161;

	wire w130161;

	wire w2020161;
	repeater #(4, 1'b1, 0, 0) c2020161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020161));
	wire w2070161;
	repeater #(2, 1'b1, 0, 0) c2070161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070161));
	wire w00162;
	repeater #(1, 1'b1, 0, 0) c00162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w00162));
	wire w20162;
	repeater #(4, 1'b1, 0, 0) c20162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20162));
	wire w70162;
	repeater #(1, 1'b0, 0, 0) c70162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70162));
	wire w100162;
	repeater #(4, 1'b0, 0, 0) c100162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100162));
	wire w150162;
	repeater #(2, 1'b1, 0, 0) c150162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150162));
	wire w2070163;
	repeater #(2, 1'b1, 0, 0) c2070163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070163));
	wire w150164;
	repeater #(2, 1'b1, 0, 0) c150164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150164));
	wire w70165;
	repeater #(1, 1'b0, 0, 0) c70165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70165));
	wire w80165;
	repeater #(1, 1'b0, 0, 0) c80165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80165));
	wire w70166;
	repeater #(4, 1'b0, 0, 0) c70166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70166));
	wire w2020166;

	wire w2030166;

	wire w2060166;
	repeater #(1, 1'b0, 0, 0) c2060166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060166));
	wire w2070166;

	wire w20167;

	wire w30167;

	wire w60167;
	repeater #(1, 1'b1, 0, 0) c60167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60167));
	wire w70167;

	wire w100167;

	wire w110167;

	wire w140167;
	repeater #(1, 1'b1, 0, 0) c140167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140167));
	wire w150167;

	wire w80169;
	torch #(1'b1) c80169 (.i_clk(tick), .i_in(), .o_out(w80169));
	wire w2020170;
	repeater #(1, 1'b1, 0, 0) c2020170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020170));
	wire w2030170;

	wire w2060170;
	repeater #(1, 1'b1, 0, 0) c2060170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2060170));
	wire w2070170;

	wire w20171;
	repeater #(1, 1'b1, 0, 0) c20171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20171));
	wire w30171;

	wire w60171;
	repeater #(1, 1'b0, 0, 0) c60171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60171));
	wire w70171;

	wire w100171;
	repeater #(1, 1'b1, 0, 0) c100171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100171));
	wire w110171;

	wire w140171;
	repeater #(1, 1'b1, 0, 0) c140171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w140171));
	wire w150171;

	wire w180171;
	repeater #(1, 1'b1, 0, 0) c180171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180171));
	wire w190171;

	wire w2020173;
	repeater #(1, 1'b1, 0, 0) c2020173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020173));
	wire w2070173;
	repeater #(1, 1'b1, 0, 0) c2070173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070173));
	wire w20174;
	repeater #(1, 1'b1, 0, 0) c20174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20174));
	wire w70174;
	repeater #(1, 1'b0, 0, 0) c70174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70174));
	wire w100174;
	repeater #(1, 1'b1, 0, 0) c100174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100174));
	wire w150174;
	repeater #(1, 1'b1, 0, 0) c150174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150174));
	wire w2040174;

	wire w2050174;

	wire w40175;

	wire w50175;

	wire w120175;

	wire w130175;

	wire w180175;
	repeater #(4, 1'b1, 0, 0) c180175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180175));
	wire w2020175;
	repeater #(4, 1'b1, 0, 0) c2020175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2020175));
	wire w2070175;
	repeater #(2, 1'b1, 0, 0) c2070175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070175));
	wire w20176;
	repeater #(4, 1'b1, 0, 0) c20176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20176));
	wire w70176;
	repeater #(2, 1'b0, 0, 0) c70176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70176));
	wire w100176;
	repeater #(4, 1'b1, 0, 0) c100176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w100176));
	wire w150176;
	repeater #(2, 1'b1, 0, 0) c150176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150176));
	wire w2070177;
	repeater #(2, 1'b1, 0, 0) c2070177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2070177));
	wire w70178;
	repeater #(2, 1'b0, 0, 0) c70178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70178));
	wire w150178;
	repeater #(2, 1'b1, 0, 0) c150178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150178));
	wire w1810;
	repeater #(2, 1'b1, 0, 0) c1810 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1810));
	wire w20211;

	wire w20311;

	wire w20611;
	repeater #(1, 1'b1, 0, 0) c20611 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20611));
	wire w20711;

	wire w212;

	wire w312;

	wire w612;
	repeater #(1, 1'b0, 0, 0) c612 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w612));
	wire w712;

	wire w1012;

	wire w1112;

	wire w1412;
	repeater #(1, 1'b1, 0, 0) c1412 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1412));
	wire w1512;

	wire w20214;
	repeater #(1, 1'b1, 0, 0) c20214 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20214));
	wire w20714;
	repeater #(1, 1'b0, 0, 0) c20714 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20714));
	wire w1015;
	repeater #(1, 1'b1, 0, 0) c1015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1015));
	wire w1515;
	repeater #(1, 1'b1, 0, 0) c1515 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1515));
	wire w20415;

	wire w20515;

	wire w116;
	repeater #(1, 1'b0, 0, 0) c116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116));
	wire w416;

	wire w516;

	wire w1216;

	wire w1316;

	wire w20216;
	repeater #(4, 1'b1, 0, 0) c20216 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20216));
	wire w20716;
	repeater #(2, 1'b0, 0, 0) c20716 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20716));
	wire w017;
	repeater #(1, 1'b0, 0, 0) c017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w017));
	wire w217;
	repeater #(4, 1'b0, 0, 0) c217 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w217));
	wire w717;
	repeater #(1, 1'b1, 0, 0) c717 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w717));
	wire w1017;
	repeater #(4, 1'b1, 0, 0) c1017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1017));
	wire w1517;
	repeater #(2, 1'b1, 0, 0) c1517 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1517));
	wire w20718;
	repeater #(2, 1'b0, 0, 0) c20718 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20718));
	wire w1519;
	repeater #(2, 1'b1, 0, 0) c1519 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1519));
	wire w7110;
	repeater #(1, 1'b1, 0, 0) c7110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7110));
	wire w8110;
	repeater #(1, 1'b1, 0, 0) c8110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8110));
	wire w7111;
	repeater #(4, 1'b1, 0, 0) c7111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7111));
	wire w202111;

	wire w203111;

	wire w206111;
	repeater #(1, 1'b0, 0, 0) c206111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206111));
	wire w207111;

	wire w2112;

	wire w3112;

	wire w6112;
	repeater #(1, 1'b1, 0, 0) c6112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6112));
	wire w7112;

	wire w10112;

	wire w11112;

	wire w14112;
	repeater #(1, 1'b1, 0, 0) c14112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14112));
	wire w15112;

	wire w8114;
	torch #(1'b0) c8114 (.i_clk(tick), .i_in(), .o_out(w8114));
	wire w202115;
	repeater #(1, 1'b1, 0, 0) c202115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202115));
	wire w203115;

	wire w206115;
	repeater #(1, 1'b1, 0, 0) c206115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206115));
	wire w207115;

	wire w2116;
	repeater #(1, 1'b1, 0, 0) c2116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2116));
	wire w3116;

	wire w6116;
	repeater #(1, 1'b0, 0, 0) c6116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6116));
	wire w7116;

	wire w10116;
	repeater #(1, 1'b1, 0, 0) c10116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10116));
	wire w11116;

	wire w14116;
	repeater #(1, 1'b1, 0, 0) c14116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14116));
	wire w15116;

	wire w18116;
	repeater #(1, 1'b1, 0, 0) c18116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18116));
	wire w19116;

	wire w202118;
	repeater #(1, 1'b1, 0, 0) c202118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202118));
	wire w207118;
	repeater #(1, 1'b1, 0, 0) c207118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207118));
	wire w2119;
	repeater #(1, 1'b1, 0, 0) c2119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2119));
	wire w7119;
	repeater #(1, 1'b0, 0, 0) c7119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7119));
	wire w10119;
	repeater #(1, 1'b1, 0, 0) c10119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10119));
	wire w15119;
	repeater #(1, 1'b1, 0, 0) c15119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15119));
	wire w204119;

	wire w205119;

	wire w4120;

	wire w5120;

	wire w12120;

	wire w13120;

	wire w18120;
	repeater #(4, 1'b1, 0, 0) c18120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18120));
	wire w202120;
	repeater #(4, 1'b1, 0, 0) c202120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202120));
	wire w207120;
	repeater #(2, 1'b1, 0, 0) c207120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207120));
	wire w2121;
	repeater #(4, 1'b1, 0, 0) c2121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2121));
	wire w7121;
	repeater #(2, 1'b0, 0, 0) c7121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7121));
	wire w10121;
	repeater #(4, 1'b1, 0, 0) c10121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10121));
	wire w15121;
	repeater #(2, 1'b1, 0, 0) c15121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15121));
	wire w207122;
	repeater #(2, 1'b1, 0, 0) c207122 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207122));
	wire w7123;
	repeater #(2, 1'b0, 0, 0) c7123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7123));
	wire w15123;
	repeater #(2, 1'b1, 0, 0) c15123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15123));
	wire w18124;
	repeater #(2, 1'b1, 0, 0) c18124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18124));
	wire w202125;

	wire w203125;

	wire w206125;
	repeater #(1, 1'b0, 0, 0) c206125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206125));
	wire w207125;

	wire w2126;

	wire w3126;

	wire w6126;
	repeater #(1, 1'b0, 0, 0) c6126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6126));
	wire w7126;

	wire w10126;

	wire w11126;

	wire w14126;
	repeater #(1, 1'b1, 0, 0) c14126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14126));
	wire w15126;

	wire w202128;
	repeater #(1, 1'b1, 0, 0) c202128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202128));
	wire w207128;
	repeater #(1, 1'b0, 0, 0) c207128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207128));
	wire w10129;
	repeater #(1, 1'b1, 0, 0) c10129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10129));
	wire w15129;
	repeater #(1, 1'b1, 0, 0) c15129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15129));
	wire w204129;

	wire w205129;

	wire w1130;
	repeater #(1, 1'b0, 0, 0) c1130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1130));
	wire w4130;

	wire w5130;

	wire w12130;

	wire w13130;

	wire w202130;
	repeater #(4, 1'b1, 0, 0) c202130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202130));
	wire w207130;
	repeater #(2, 1'b0, 0, 0) c207130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207130));
	wire w0131;
	repeater #(1, 1'b0, 0, 0) c0131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0131));
	wire w2131;
	repeater #(4, 1'b0, 0, 0) c2131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2131));
	wire w7131;
	repeater #(1, 1'b1, 0, 0) c7131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7131));
	wire w10131;
	repeater #(4, 1'b1, 0, 0) c10131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10131));
	wire w15131;
	repeater #(2, 1'b1, 0, 0) c15131 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15131));
	wire w207132;
	repeater #(2, 1'b0, 0, 0) c207132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207132));
	wire w15133;
	repeater #(2, 1'b1, 0, 0) c15133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15133));
	wire w7134;
	repeater #(1, 1'b1, 0, 0) c7134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7134));
	wire w8134;
	repeater #(1, 1'b1, 0, 0) c8134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8134));
	wire w7135;
	repeater #(4, 1'b1, 0, 0) c7135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7135));
	wire w202135;

	wire w203135;

	wire w206135;
	repeater #(1, 1'b0, 0, 0) c206135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206135));
	wire w207135;

	wire w2136;

	wire w3136;

	wire w6136;
	repeater #(1, 1'b1, 0, 0) c6136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6136));
	wire w7136;

	wire w10136;

	wire w11136;

	wire w14136;
	repeater #(1, 1'b1, 0, 0) c14136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14136));
	wire w15136;

	wire w8138;
	torch #(1'b0) c8138 (.i_clk(tick), .i_in(), .o_out(w8138));
	wire w202139;
	repeater #(1, 1'b0, 0, 0) c202139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202139));
	wire w203139;

	wire w206139;
	repeater #(1, 1'b0, 0, 0) c206139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206139));
	wire w207139;

	wire w2140;
	repeater #(1, 1'b0, 0, 0) c2140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2140));
	wire w3140;

	wire w6140;
	repeater #(1, 1'b0, 0, 0) c6140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6140));
	wire w7140;

	wire w10140;
	repeater #(1, 1'b0, 0, 0) c10140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10140));
	wire w11140;

	wire w14140;
	repeater #(1, 1'b0, 0, 0) c14140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14140));
	wire w15140;

	wire w18140;
	repeater #(1, 1'b0, 0, 0) c18140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18140));
	wire w19140;

	wire w202142;
	repeater #(1, 1'b0, 0, 0) c202142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202142));
	wire w207142;
	repeater #(1, 1'b0, 0, 0) c207142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207142));
	wire w2143;
	repeater #(1, 1'b0, 0, 0) c2143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2143));
	wire w7143;
	repeater #(1, 1'b0, 0, 0) c7143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7143));
	wire w10143;
	repeater #(1, 1'b0, 0, 0) c10143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10143));
	wire w15143;
	repeater #(1, 1'b0, 0, 0) c15143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15143));
	wire w204143;

	wire w205143;

	wire w4144;

	wire w5144;

	wire w12144;

	wire w13144;

	wire w18144;
	repeater #(4, 1'b0, 0, 0) c18144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18144));
	wire w202144;
	repeater #(4, 1'b0, 0, 0) c202144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202144));
	wire w207144;
	repeater #(2, 1'b0, 0, 0) c207144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207144));
	wire w2145;
	repeater #(4, 1'b0, 0, 0) c2145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2145));
	wire w7145;
	repeater #(2, 1'b0, 0, 0) c7145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7145));
	wire w10145;
	repeater #(4, 1'b0, 0, 0) c10145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10145));
	wire w15145;
	repeater #(2, 1'b0, 0, 0) c15145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15145));
	wire w207146;
	repeater #(2, 1'b0, 0, 0) c207146 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207146));
	wire w7147;
	repeater #(2, 1'b0, 0, 0) c7147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7147));
	wire w15147;
	repeater #(2, 1'b0, 0, 0) c15147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15147));
	wire w18148;
	repeater #(2, 1'b0, 0, 0) c18148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18148));
	wire w202149;

	wire w203149;

	wire w206149;
	repeater #(1, 1'b0, 0, 0) c206149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206149));
	wire w207149;

	wire w2150;

	wire w3150;

	wire w6150;
	repeater #(1, 1'b0, 0, 0) c6150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6150));
	wire w7150;

	wire w10150;

	wire w11150;

	wire w14150;
	repeater #(1, 1'b0, 0, 0) c14150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14150));
	wire w15150;

	wire w202152;
	repeater #(1, 1'b0, 0, 0) c202152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202152));
	wire w207152;
	repeater #(1, 1'b0, 0, 0) c207152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207152));
	wire w10153;
	repeater #(1, 1'b0, 0, 0) c10153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10153));
	wire w15153;
	repeater #(1, 1'b0, 0, 0) c15153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15153));
	wire w204153;

	wire w205153;

	wire w1154;
	repeater #(1, 1'b0, 0, 0) c1154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1154));
	wire w4154;

	wire w5154;

	wire w12154;

	wire w13154;

	wire w202154;
	repeater #(4, 1'b0, 0, 0) c202154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202154));
	wire w207154;
	repeater #(2, 1'b0, 0, 0) c207154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207154));
	wire w0155;
	repeater #(1, 1'b0, 0, 0) c0155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0155));
	wire w2155;
	repeater #(4, 1'b0, 0, 0) c2155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2155));
	wire w7155;
	repeater #(1, 1'b0, 0, 0) c7155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7155));
	wire w10155;
	repeater #(4, 1'b0, 0, 0) c10155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10155));
	wire w15155;
	repeater #(2, 1'b0, 0, 0) c15155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15155));
	wire w207156;
	repeater #(2, 1'b0, 0, 0) c207156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207156));
	wire w15157;
	repeater #(2, 1'b0, 0, 0) c15157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15157));
	wire w7158;
	repeater #(1, 1'b0, 0, 0) c7158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7158));
	wire w8158;
	repeater #(1, 1'b0, 0, 0) c8158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8158));
	wire w7159;
	repeater #(4, 1'b0, 0, 0) c7159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7159));
	wire w202159;

	wire w203159;

	wire w206159;
	repeater #(1, 1'b0, 0, 0) c206159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206159));
	wire w207159;

	wire w2160;

	wire w3160;

	wire w6160;
	repeater #(1, 1'b0, 0, 0) c6160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6160));
	wire w7160;

	wire w10160;

	wire w11160;

	wire w14160;
	repeater #(1, 1'b0, 0, 0) c14160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14160));
	wire w15160;

	wire w8162;
	torch #(1'b0) c8162 (.i_clk(tick), .i_in(), .o_out(w8162));
	wire w202163;
	repeater #(1, 1'b1, 0, 0) c202163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202163));
	wire w203163;

	wire w206163;
	repeater #(1, 1'b1, 0, 0) c206163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206163));
	wire w207163;

	wire w2164;
	repeater #(1, 1'b1, 0, 0) c2164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2164));
	wire w3164;

	wire w6164;
	repeater #(1, 1'b1, 0, 0) c6164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6164));
	wire w7164;

	wire w10164;
	repeater #(1, 1'b1, 0, 0) c10164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10164));
	wire w11164;

	wire w14164;
	repeater #(1, 1'b1, 0, 0) c14164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14164));
	wire w15164;

	wire w18164;
	repeater #(1, 1'b1, 0, 0) c18164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18164));
	wire w19164;

	wire w202166;
	repeater #(1, 1'b1, 0, 0) c202166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202166));
	wire w207166;
	repeater #(1, 1'b1, 0, 0) c207166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207166));
	wire w2167;
	repeater #(1, 1'b1, 0, 0) c2167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2167));
	wire w7167;
	repeater #(1, 1'b1, 0, 0) c7167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7167));
	wire w10167;
	repeater #(1, 1'b1, 0, 0) c10167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10167));
	wire w15167;
	repeater #(1, 1'b1, 0, 0) c15167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15167));
	wire w204167;

	wire w205167;

	wire w4168;

	wire w5168;

	wire w12168;

	wire w13168;

	wire w18168;
	repeater #(4, 1'b1, 0, 0) c18168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18168));
	wire w202168;
	repeater #(4, 1'b1, 0, 0) c202168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202168));
	wire w207168;
	repeater #(2, 1'b1, 0, 0) c207168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207168));
	wire w2169;
	repeater #(4, 1'b1, 0, 0) c2169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2169));
	wire w7169;
	repeater #(2, 1'b1, 0, 0) c7169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7169));
	wire w10169;
	repeater #(4, 1'b1, 0, 0) c10169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10169));
	wire w15169;
	repeater #(2, 1'b1, 0, 0) c15169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15169));
	wire w207170;
	repeater #(2, 1'b1, 0, 0) c207170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207170));
	wire w7171;
	repeater #(2, 1'b1, 0, 0) c7171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7171));
	wire w15171;
	repeater #(2, 1'b1, 0, 0) c15171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15171));
	wire w18172;
	repeater #(2, 1'b1, 0, 0) c18172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18172));
	wire w202173;

	wire w203173;

	wire w206173;
	repeater #(1, 1'b0, 0, 0) c206173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206173));
	wire w207173;

	wire w2174;

	wire w3174;

	wire w6174;
	repeater #(1, 1'b0, 0, 0) c6174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6174));
	wire w7174;

	wire w10174;

	wire w11174;

	wire w14174;
	repeater #(1, 1'b0, 0, 0) c14174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14174));
	wire w15174;

	wire w202176;
	repeater #(1, 1'b1, 0, 0) c202176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202176));
	wire w207176;
	repeater #(1, 1'b1, 0, 0) c207176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207176));
	wire w10177;
	repeater #(1, 1'b1, 0, 0) c10177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10177));
	wire w15177;
	repeater #(1, 1'b1, 0, 0) c15177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15177));
	wire w204177;

	wire w205177;

	wire w1178;
	repeater #(1, 1'b1, 0, 0) c1178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1178));
	wire w4178;

	wire w5178;

	wire w12178;

	wire w13178;

	wire w202178;
	repeater #(4, 1'b1, 0, 0) c202178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202178));
	wire w207178;
	repeater #(2, 1'b1, 0, 0) c207178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207178));
	wire w0179;
	repeater #(1, 1'b1, 0, 0) c0179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w0179));
	wire w2179;
	repeater #(4, 1'b1, 0, 0) c2179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2179));
	wire w7179;
	repeater #(1, 1'b1, 0, 0) c7179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7179));
	wire w10179;
	repeater #(4, 1'b1, 0, 0) c10179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10179));
	wire w15179;
	repeater #(2, 1'b1, 0, 0) c15179 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15179));
	wire w207180;
	repeater #(2, 1'b1, 0, 0) c207180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207180));
	wire w15181;
	repeater #(2, 1'b1, 0, 0) c15181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15181));
	wire w7182;
	repeater #(1, 1'b1, 0, 0) c7182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7182));
	wire w8182;
	repeater #(1, 1'b1, 0, 0) c8182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8182));
	wire w7183;
	repeater #(4, 1'b1, 0, 0) c7183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w7183));
	wire w202183;

	wire w203183;

	wire w206183;
	repeater #(1, 1'b0, 0, 0) c206183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206183));
	wire w207183;

	wire w2184;

	wire w3184;

	wire w6184;
	repeater #(1, 1'b0, 0, 0) c6184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6184));
	wire w7184;

	wire w10184;

	wire w11184;

	wire w14184;
	repeater #(1, 1'b1, 0, 0) c14184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14184));
	wire w15184;

	wire w8186;
	torch #(1'b1) c8186 (.i_clk(tick), .i_in(), .o_out(w8186));
	wire w18503;
	repeater #(1, 1'b0, 0, 0) c18503 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18503));
	wire w18604;
	repeater #(1, 1'b0, 0, 0) c18604 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18604));
	wire w14805;
	repeater #(1, 1'b0, 0, 0) c14805 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14805));
	wire w16505;
	repeater #(2, 1'b0, 0, 0) c16505 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16505));
	wire w16605;
	repeater #(1, 1'b0, 0, 0) c16605 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16605));
	wire w16705;

	wire w18205;

	wire w18505;
	repeater #(1, 1'b0, 0, 0) c18505 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18505));
	wire w19505;
	repeater #(1, 1'b0, 0, 0) c19505 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19505));
	wire w20005;
	repeater #(1, 1'b1, 0, 0) c20005 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w20005));
	wire w18406;
	repeater #(1, 1'b0, 0, 0) c18406 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18406));
	wire w19706;

	wire w19806;

	wire w19808;
	repeater #(1, 1'b1, 0, 0) c19808 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w19808));
	wire w409;
	repeater #(1, 1'b1, 0, 0) c409 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w409));
	wire w4010;

	wire w6011;
	repeater #(1, 1'b0, 0, 0) c6011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6011));
	wire w183011;
	repeater #(1, 1'b0, 0, 0) c183011 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183011));
	wire w145019;
	repeater #(1, 1'b1, 0, 0) c145019 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w145019));
	wire w6027;
	repeater #(1, 1'b0, 0, 0) c6027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6027));
	wire w4033;
	repeater #(1, 1'b1, 0, 0) c4033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4033));
	wire w4034;

	wire w6035;
	repeater #(1, 1'b0, 0, 0) c6035 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6035));
	wire w6051;
	repeater #(1, 1'b0, 0, 0) c6051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6051));
	wire w4057;
	repeater #(1, 1'b1, 0, 0) c4057 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4057));
	wire w4058;

	wire w6059;
	repeater #(1, 1'b0, 0, 0) c6059 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6059));
	wire w6075;
	repeater #(1, 1'b0, 0, 0) c6075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6075));
	wire w4081;
	repeater #(1, 1'b1, 0, 0) c4081 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w4081));
	wire w4082;

	wire w6083;
	repeater #(1, 1'b0, 0, 0) c6083 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6083));
	wire w6099;
	repeater #(1, 1'b0, 0, 0) c6099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w6099));
	wire w40105;
	repeater #(1, 1'b1, 0, 0) c40105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w40105));
	wire w40106;

	wire w60107;
	repeater #(1, 1'b0, 0, 0) c60107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60107));
	wire w60123;
	repeater #(1, 1'b0, 0, 0) c60123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w60123));
	wire w80128;
	repeater #(1, 1'b0, 0, 0) c80128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w80128));
	wire w90130;

	wire w120130;
	assign outputs[122] = ();
	wire w90131;

	wire w70132;
	repeater #(1, 1'b0, 0, 0) c70132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w70132));
	wire w14915;

	wire w186110;
	repeater #(1, 1'b1, 0, 0) c186110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186110));
	wire w187110;

	wire w190110;
	repeater #(1, 1'b1, 0, 0) c190110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190110));
	wire w191110;

	wire w194110;
	repeater #(1, 1'b1, 0, 0) c194110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194110));
	wire w195110;

	wire w198110;
	repeater #(1, 1'b1, 0, 0) c198110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198110));
	wire w199110;

	wire w202110;
	repeater #(1, 1'b1, 0, 0) c202110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202110));
	wire w203110;

	wire w206110;
	repeater #(1, 1'b0, 0, 0) c206110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206110));
	wire w207110;

	wire w2111;
	repeater #(1, 1'b0, 0, 0) c2111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2111));
	wire w3111;

	wire w186113;
	repeater #(1, 1'b1, 0, 0) c186113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186113));
	wire w191113;
	repeater #(1, 1'b1, 0, 0) c191113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191113));
	wire w194113;
	repeater #(1, 1'b1, 0, 0) c194113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194113));
	wire w199113;
	repeater #(1, 1'b1, 0, 0) c199113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199113));
	wire w202113;
	repeater #(1, 1'b1, 0, 0) c202113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202113));
	wire w207113;
	repeater #(1, 1'b0, 0, 0) c207113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207113));
	wire w188114;

	wire w189114;

	wire w196114;

	wire w197114;

	wire w204114;

	wire w205114;

	wire w2115;
	repeater #(4, 1'b0, 0, 0) c2115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2115));
	wire w186115;
	repeater #(4, 1'b1, 0, 0) c186115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186115));
	wire w191115;
	repeater #(2, 1'b1, 0, 0) c191115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191115));
	wire w194115;
	repeater #(4, 1'b1, 0, 0) c194115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194115));
	wire w199115;
	repeater #(2, 1'b1, 0, 0) c199115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199115));
	wire w202115;
	repeater #(4, 1'b1, 0, 0) c202115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202115));
	wire w207115;
	repeater #(2, 1'b0, 0, 0) c207115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207115));
	wire w191117;
	repeater #(2, 1'b1, 0, 0) c191117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191117));
	wire w199117;
	repeater #(2, 1'b1, 0, 0) c199117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199117));
	wire w207117;
	repeater #(2, 1'b0, 0, 0) c207117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207117));
	wire w146118;

	wire w2119;
	repeater #(2, 1'b0, 0, 0) c2119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2119));
	wire w186120;

	wire w187120;

	wire w190120;
	repeater #(1, 1'b0, 0, 0) c190120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190120));
	wire w191120;

	wire w194120;

	wire w195120;

	wire w198120;
	repeater #(1, 1'b1, 0, 0) c198120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198120));
	wire w199120;

	wire w202120;

	wire w203120;

	wire w206120;
	repeater #(1, 1'b1, 0, 0) c206120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206120));
	wire w207120;

	wire w186123;
	repeater #(1, 1'b1, 0, 0) c186123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186123));
	wire w191123;
	repeater #(1, 1'b1, 0, 0) c191123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191123));
	wire w202123;
	repeater #(1, 1'b1, 0, 0) c202123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202123));
	wire w207123;
	repeater #(1, 1'b0, 0, 0) c207123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207123));
	wire w188124;

	wire w189124;

	wire w193124;
	repeater #(1, 1'b1, 0, 0) c193124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193124));
	wire w196124;

	wire w197124;

	wire w204124;

	wire w205124;

	wire w186125;
	repeater #(4, 1'b1, 0, 0) c186125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186125));
	wire w191125;
	repeater #(2, 1'b1, 0, 0) c191125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191125));
	wire w192125;
	repeater #(1, 1'b1, 0, 0) c192125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192125));
	wire w194125;
	repeater #(4, 1'b1, 0, 0) c194125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194125));
	wire w199125;
	repeater #(1, 1'b1, 0, 0) c199125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199125));
	wire w202125;
	repeater #(4, 1'b1, 0, 0) c202125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202125));
	wire w207125;
	repeater #(2, 1'b0, 0, 0) c207125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207125));
	wire w191127;
	repeater #(2, 1'b1, 0, 0) c191127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191127));
	wire w207127;
	repeater #(2, 1'b0, 0, 0) c207127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207127));
	wire w199128;
	repeater #(1, 1'b1, 0, 0) c199128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199128));
	wire w200128;
	repeater #(1, 1'b1, 0, 0) c200128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200128));
	wire w199129;
	repeater #(4, 1'b1, 0, 0) c199129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199129));
	wire w186130;

	wire w187130;

	wire w190130;
	repeater #(1, 1'b0, 0, 0) c190130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190130));
	wire w191130;

	wire w194130;

	wire w195130;

	wire w198130;
	repeater #(1, 1'b1, 0, 0) c198130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198130));
	wire w199130;

	wire w202130;

	wire w203130;

	wire w206130;
	repeater #(1, 1'b1, 0, 0) c206130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206130));
	wire w207130;

	wire w200132;
	torch #(1'b1) c200132 (.i_clk(tick), .i_in(), .o_out(w200132));
	wire w186134;
	repeater #(1, 1'b0, 0, 0) c186134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186134));
	wire w187134;

	wire w190134;
	repeater #(1, 1'b0, 0, 0) c190134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190134));
	wire w191134;

	wire w194134;
	repeater #(1, 1'b0, 0, 0) c194134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194134));
	wire w195134;

	wire w198134;
	repeater #(1, 1'b1, 0, 0) c198134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198134));
	wire w199134;

	wire w202134;
	repeater #(1, 1'b0, 0, 0) c202134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202134));
	wire w203134;

	wire w206134;
	repeater #(1, 1'b0, 0, 0) c206134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206134));
	wire w207134;

	wire w2135;
	repeater #(1, 1'b0, 0, 0) c2135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2135));
	wire w3135;

	wire w186137;
	repeater #(1, 1'b0, 0, 0) c186137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186137));
	wire w191137;
	repeater #(1, 1'b0, 0, 0) c191137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191137));
	wire w194137;
	repeater #(1, 1'b0, 0, 0) c194137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194137));
	wire w199137;
	repeater #(1, 1'b1, 0, 0) c199137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199137));
	wire w202137;
	repeater #(1, 1'b0, 0, 0) c202137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202137));
	wire w207137;
	repeater #(1, 1'b0, 0, 0) c207137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207137));
	wire w188138;

	wire w189138;

	wire w196138;

	wire w197138;

	wire w204138;

	wire w205138;

	wire w2139;
	repeater #(4, 1'b0, 0, 0) c2139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2139));
	wire w186139;
	repeater #(4, 1'b0, 0, 0) c186139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186139));
	wire w191139;
	repeater #(2, 1'b0, 0, 0) c191139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191139));
	wire w194139;
	repeater #(4, 1'b0, 0, 0) c194139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194139));
	wire w199139;
	repeater #(2, 1'b1, 0, 0) c199139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199139));
	wire w202139;
	repeater #(4, 1'b0, 0, 0) c202139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202139));
	wire w207139;
	repeater #(2, 1'b0, 0, 0) c207139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207139));
	wire w191141;
	repeater #(2, 1'b0, 0, 0) c191141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191141));
	wire w199141;
	repeater #(2, 1'b1, 0, 0) c199141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199141));
	wire w207141;
	repeater #(2, 1'b0, 0, 0) c207141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207141));
	wire w2143;
	repeater #(2, 1'b0, 0, 0) c2143 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2143));
	wire w186144;

	wire w187144;

	wire w190144;
	repeater #(1, 1'b1, 0, 0) c190144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190144));
	wire w191144;

	wire w194144;

	wire w195144;

	wire w198144;
	repeater #(1, 1'b0, 0, 0) c198144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198144));
	wire w199144;

	wire w202144;

	wire w203144;

	wire w206144;
	repeater #(1, 1'b1, 0, 0) c206144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206144));
	wire w207144;

	wire w186147;
	repeater #(1, 1'b0, 0, 0) c186147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186147));
	wire w191147;
	repeater #(1, 1'b1, 0, 0) c191147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191147));
	wire w202147;
	repeater #(1, 1'b0, 0, 0) c202147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202147));
	wire w207147;
	repeater #(1, 1'b0, 0, 0) c207147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207147));
	wire w188148;

	wire w189148;

	wire w193148;
	repeater #(1, 1'b1, 0, 0) c193148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193148));
	wire w196148;

	wire w197148;

	wire w204148;

	wire w205148;

	wire w186149;
	repeater #(4, 1'b0, 0, 0) c186149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186149));
	wire w191149;
	repeater #(2, 1'b1, 0, 0) c191149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191149));
	wire w192149;
	repeater #(1, 1'b1, 0, 0) c192149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192149));
	wire w194149;
	repeater #(4, 1'b1, 0, 0) c194149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194149));
	wire w199149;
	repeater #(1, 1'b0, 0, 0) c199149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199149));
	wire w202149;
	repeater #(4, 1'b0, 0, 0) c202149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202149));
	wire w207149;
	repeater #(2, 1'b0, 0, 0) c207149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207149));
	wire w191151;
	repeater #(2, 1'b1, 0, 0) c191151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191151));
	wire w207151;
	repeater #(2, 1'b0, 0, 0) c207151 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207151));
	wire w199152;
	repeater #(1, 1'b0, 0, 0) c199152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199152));
	wire w200152;
	repeater #(1, 1'b0, 0, 0) c200152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200152));
	wire w199153;
	repeater #(4, 1'b0, 0, 0) c199153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199153));
	wire w186154;

	wire w187154;

	wire w190154;
	repeater #(1, 1'b0, 0, 0) c190154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190154));
	wire w191154;

	wire w194154;

	wire w195154;

	wire w198154;
	repeater #(1, 1'b1, 0, 0) c198154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198154));
	wire w199154;

	wire w202154;

	wire w203154;

	wire w206154;
	repeater #(1, 1'b1, 0, 0) c206154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206154));
	wire w207154;

	wire w200156;
	torch #(1'b1) c200156 (.i_clk(tick), .i_in(), .o_out(w200156));
	wire w186158;
	repeater #(1, 1'b0, 0, 0) c186158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186158));
	wire w187158;

	wire w190158;
	repeater #(1, 1'b0, 0, 0) c190158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190158));
	wire w191158;

	wire w194158;
	repeater #(1, 1'b0, 0, 0) c194158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194158));
	wire w195158;

	wire w198158;
	repeater #(1, 1'b1, 0, 0) c198158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198158));
	wire w199158;

	wire w202158;
	repeater #(1, 1'b0, 0, 0) c202158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202158));
	wire w203158;

	wire w206158;
	repeater #(1, 1'b1, 0, 0) c206158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206158));
	wire w207158;

	wire w2159;
	repeater #(1, 1'b1, 0, 0) c2159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2159));
	wire w3159;

	wire w186161;
	repeater #(1, 1'b0, 0, 0) c186161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186161));
	wire w191161;
	repeater #(1, 1'b0, 0, 0) c191161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191161));
	wire w194161;
	repeater #(1, 1'b0, 0, 0) c194161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194161));
	wire w199161;
	repeater #(1, 1'b1, 0, 0) c199161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199161));
	wire w202161;
	repeater #(1, 1'b0, 0, 0) c202161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202161));
	wire w207161;
	repeater #(1, 1'b1, 0, 0) c207161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207161));
	wire w188162;

	wire w189162;

	wire w196162;

	wire w197162;

	wire w204162;

	wire w205162;

	wire w2163;
	repeater #(4, 1'b1, 0, 0) c2163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2163));
	wire w186163;
	repeater #(4, 1'b0, 0, 0) c186163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186163));
	wire w191163;
	repeater #(2, 1'b0, 0, 0) c191163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191163));
	wire w194163;
	repeater #(4, 1'b0, 0, 0) c194163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194163));
	wire w199163;
	repeater #(2, 1'b1, 0, 0) c199163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199163));
	wire w202163;
	repeater #(4, 1'b0, 0, 0) c202163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202163));
	wire w207163;
	repeater #(2, 1'b1, 0, 0) c207163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207163));
	wire w191165;
	repeater #(2, 1'b0, 0, 0) c191165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191165));
	wire w199165;
	repeater #(2, 1'b1, 0, 0) c199165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199165));
	wire w207165;
	repeater #(2, 1'b1, 0, 0) c207165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207165));
	wire w2167;
	repeater #(2, 1'b1, 0, 0) c2167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2167));
	wire w186168;

	wire w187168;

	wire w190168;
	repeater #(1, 1'b0, 0, 0) c190168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190168));
	wire w191168;

	wire w194168;

	wire w195168;

	wire w198168;
	repeater #(1, 1'b0, 0, 0) c198168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198168));
	wire w199168;

	wire w202168;

	wire w203168;

	wire w206168;
	repeater #(1, 1'b1, 0, 0) c206168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206168));
	wire w207168;

	wire w186171;
	repeater #(1, 1'b0, 0, 0) c186171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186171));
	wire w191171;
	repeater #(1, 1'b1, 0, 0) c191171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191171));
	wire w202171;
	repeater #(1, 1'b0, 0, 0) c202171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202171));
	wire w207171;
	repeater #(1, 1'b1, 0, 0) c207171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207171));
	wire w188172;

	wire w189172;

	wire w193172;
	repeater #(1, 1'b1, 0, 0) c193172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193172));
	wire w196172;

	wire w197172;

	wire w204172;

	wire w205172;

	wire w186173;
	repeater #(4, 1'b0, 0, 0) c186173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186173));
	wire w191173;
	repeater #(2, 1'b1, 0, 0) c191173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191173));
	wire w192173;
	repeater #(1, 1'b1, 0, 0) c192173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192173));
	wire w194173;
	repeater #(4, 1'b1, 0, 0) c194173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194173));
	wire w199173;
	repeater #(1, 1'b0, 0, 0) c199173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199173));
	wire w202173;
	repeater #(4, 1'b0, 0, 0) c202173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202173));
	wire w207173;
	repeater #(2, 1'b1, 0, 0) c207173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207173));
	wire w191175;
	repeater #(2, 1'b1, 0, 0) c191175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191175));
	wire w207175;
	repeater #(2, 1'b1, 0, 0) c207175 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207175));
	wire w199176;
	repeater #(1, 1'b0, 0, 0) c199176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199176));
	wire w200176;
	repeater #(1, 1'b0, 0, 0) c200176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w200176));
	wire w199177;
	repeater #(4, 1'b0, 0, 0) c199177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199177));
	wire w186178;

	wire w187178;

	wire w190178;
	repeater #(1, 1'b0, 0, 0) c190178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190178));
	wire w191178;

	wire w194178;

	wire w195178;

	wire w198178;
	repeater #(1, 1'b1, 0, 0) c198178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198178));
	wire w199178;

	wire w202178;

	wire w203178;

	wire w206178;
	repeater #(1, 1'b1, 0, 0) c206178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206178));
	wire w207178;

	wire w200180;
	torch #(1'b1) c200180 (.i_clk(tick), .i_in(), .o_out(w200180));
	wire w186182;
	repeater #(1, 1'b0, 0, 0) c186182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186182));
	wire w187182;

	wire w190182;
	repeater #(1, 1'b0, 0, 0) c190182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190182));
	wire w191182;

	wire w194182;
	repeater #(1, 1'b0, 0, 0) c194182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194182));
	wire w195182;

	wire w198182;
	repeater #(1, 1'b0, 0, 0) c198182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198182));
	wire w199182;

	wire w202182;
	repeater #(1, 1'b0, 0, 0) c202182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202182));
	wire w203182;

	wire w206182;
	repeater #(1, 1'b0, 0, 0) c206182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206182));
	wire w207182;

	wire w2183;
	repeater #(1, 1'b0, 0, 0) c2183 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2183));
	wire w3183;

	wire w186185;
	repeater #(1, 1'b0, 0, 0) c186185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186185));
	wire w191185;
	repeater #(1, 1'b0, 0, 0) c191185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191185));
	wire w194185;
	repeater #(1, 1'b0, 0, 0) c194185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194185));
	wire w199185;
	repeater #(1, 1'b0, 0, 0) c199185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199185));
	wire w202185;
	repeater #(1, 1'b0, 0, 0) c202185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202185));
	wire w207185;
	repeater #(1, 1'b0, 0, 0) c207185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207185));
	wire w188186;

	wire w189186;

	wire w196186;

	wire w197186;

	wire w204186;

	wire w205186;

	wire w2187;
	repeater #(4, 1'b0, 0, 0) c2187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2187));
	wire w186187;
	repeater #(4, 1'b0, 0, 0) c186187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186187));
	wire w191187;
	repeater #(2, 1'b0, 0, 0) c191187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191187));
	wire w194187;
	repeater #(4, 1'b0, 0, 0) c194187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194187));
	wire w199187;
	repeater #(2, 1'b0, 0, 0) c199187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199187));
	wire w202187;
	repeater #(4, 1'b0, 0, 0) c202187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202187));
	wire w207187;
	repeater #(2, 1'b0, 0, 0) c207187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207187));
	wire w191189;
	repeater #(2, 1'b0, 0, 0) c191189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191189));
	wire w199189;
	repeater #(2, 1'b0, 0, 0) c199189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199189));
	wire w207189;
	repeater #(2, 1'b0, 0, 0) c207189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207189));
	wire w2191;
	repeater #(2, 1'b0, 0, 0) c2191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2191));
	wire w186192;

	wire w187192;

	wire w190192;
	repeater #(1, 1'b0, 0, 0) c190192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190192));
	wire w191192;

	wire w194192;

	wire w195192;

	wire w198192;
	repeater #(1, 1'b0, 0, 0) c198192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198192));
	wire w199192;

	wire w202192;

	wire w203192;

	wire w206192;
	repeater #(1, 1'b0, 0, 0) c206192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w206192));
	wire w207192;

	wire w186195;
	repeater #(1, 1'b0, 0, 0) c186195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186195));
	wire w191195;
	repeater #(1, 1'b0, 0, 0) c191195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191195));
	wire w202195;
	repeater #(1, 1'b0, 0, 0) c202195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202195));
	wire w207195;
	repeater #(1, 1'b0, 0, 0) c207195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207195));
	wire w188196;

	wire w189196;

	wire w193196;
	repeater #(1, 1'b0, 0, 0) c193196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w193196));
	wire w196196;

	wire w197196;

	wire w204196;

	wire w205196;

	wire w186197;
	repeater #(4, 1'b0, 0, 0) c186197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186197));
	wire w191197;
	repeater #(2, 1'b0, 0, 0) c191197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191197));
	wire w192197;
	repeater #(1, 1'b0, 0, 0) c192197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w192197));
	wire w194197;
	repeater #(4, 1'b0, 0, 0) c194197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194197));
	wire w199197;
	repeater #(1, 1'b0, 0, 0) c199197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w199197));
	wire w202197;
	repeater #(4, 1'b0, 0, 0) c202197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w202197));
	wire w207197;
	repeater #(2, 1'b0, 0, 0) c207197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207197));
	wire w191199;
	repeater #(2, 1'b0, 0, 0) c191199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191199));
	wire w207199;
	repeater #(2, 1'b0, 0, 0) c207199 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w207199));
	wire w1991100;
	repeater #(1, 1'b0, 0, 0) c1991100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991100));
	wire w2001100;
	repeater #(1, 1'b0, 0, 0) c2001100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2001100));
	wire w1991101;
	repeater #(4, 1'b0, 0, 0) c1991101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991101));
	wire w1861102;

	wire w1871102;

	wire w1901102;
	repeater #(1, 1'b0, 0, 0) c1901102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901102));
	wire w1911102;

	wire w1941102;

	wire w1951102;

	wire w1981102;
	repeater #(1, 1'b0, 0, 0) c1981102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1981102));
	wire w1991102;

	wire w2021102;

	wire w2031102;

	wire w2061102;
	repeater #(1, 1'b0, 0, 0) c2061102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2061102));
	wire w2071102;

	wire w2001104;
	torch #(1'b0) c2001104 (.i_clk(tick), .i_in(), .o_out(w2001104));
	wire w1861106;
	repeater #(1, 1'b1, 0, 0) c1861106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861106));
	wire w1871106;

	wire w1901106;
	repeater #(1, 1'b1, 0, 0) c1901106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901106));
	wire w1911106;

	wire w1941106;
	repeater #(1, 1'b1, 0, 0) c1941106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941106));
	wire w1951106;

	wire w1981106;
	repeater #(1, 1'b1, 0, 0) c1981106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1981106));
	wire w1991106;

	wire w2021106;
	repeater #(1, 1'b1, 0, 0) c2021106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021106));
	wire w2031106;

	wire w2061106;
	repeater #(1, 1'b1, 0, 0) c2061106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2061106));
	wire w2071106;

	wire w21107;
	repeater #(1, 1'b0, 0, 0) c21107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21107));
	wire w31107;

	wire w1861109;
	repeater #(1, 1'b1, 0, 0) c1861109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861109));
	wire w1911109;
	repeater #(1, 1'b1, 0, 0) c1911109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911109));
	wire w1941109;
	repeater #(1, 1'b1, 0, 0) c1941109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941109));
	wire w1991109;
	repeater #(1, 1'b1, 0, 0) c1991109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991109));
	wire w2021109;
	repeater #(1, 1'b1, 0, 0) c2021109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021109));
	wire w2071109;
	repeater #(1, 1'b1, 0, 0) c2071109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071109));
	wire w1881110;

	wire w1891110;

	wire w1961110;

	wire w1971110;

	wire w2041110;

	wire w2051110;

	wire w21111;
	repeater #(4, 1'b0, 0, 0) c21111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21111));
	wire w1861111;
	repeater #(4, 1'b1, 0, 0) c1861111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861111));
	wire w1911111;
	repeater #(2, 1'b1, 0, 0) c1911111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911111));
	wire w1941111;
	repeater #(4, 1'b1, 0, 0) c1941111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941111));
	wire w1991111;
	repeater #(2, 1'b1, 0, 0) c1991111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991111));
	wire w2021111;
	repeater #(4, 1'b1, 0, 0) c2021111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021111));
	wire w2071111;
	repeater #(2, 1'b1, 0, 0) c2071111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071111));
	wire w1911113;
	repeater #(2, 1'b1, 0, 0) c1911113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911113));
	wire w1991113;
	repeater #(2, 1'b1, 0, 0) c1991113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991113));
	wire w2071113;
	repeater #(2, 1'b1, 0, 0) c2071113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071113));
	wire w21115;
	repeater #(2, 1'b0, 0, 0) c21115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w21115));
	wire w1861116;

	wire w1871116;

	wire w1901116;
	repeater #(1, 1'b0, 0, 0) c1901116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901116));
	wire w1911116;

	wire w1941116;

	wire w1951116;

	wire w1981116;
	repeater #(1, 1'b0, 0, 0) c1981116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1981116));
	wire w1991116;

	wire w2021116;

	wire w2031116;

	wire w2061116;
	repeater #(1, 1'b0, 0, 0) c2061116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2061116));
	wire w2071116;

	wire w1861119;
	repeater #(1, 1'b1, 0, 0) c1861119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861119));
	wire w1911119;
	repeater #(1, 1'b1, 0, 0) c1911119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911119));
	wire w2021119;
	repeater #(1, 1'b1, 0, 0) c2021119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021119));
	wire w2071119;
	repeater #(1, 1'b0, 0, 0) c2071119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071119));
	wire w1881120;

	wire w1891120;

	wire w1931120;
	repeater #(1, 1'b1, 0, 0) c1931120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1931120));
	wire w1961120;

	wire w1971120;

	wire w2041120;

	wire w2051120;

	wire w1861121;
	repeater #(4, 1'b1, 0, 0) c1861121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861121));
	wire w1911121;
	repeater #(2, 1'b1, 0, 0) c1911121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911121));
	wire w1921121;
	repeater #(1, 1'b1, 0, 0) c1921121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1921121));
	wire w1941121;
	repeater #(4, 1'b1, 0, 0) c1941121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941121));
	wire w1991121;
	repeater #(1, 1'b1, 0, 0) c1991121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991121));
	wire w2021121;
	repeater #(4, 1'b1, 0, 0) c2021121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2021121));
	wire w2071121;
	repeater #(2, 1'b0, 0, 0) c2071121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071121));
	wire w1911123;
	repeater #(2, 1'b1, 0, 0) c1911123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911123));
	wire w2071123;
	repeater #(2, 1'b0, 0, 0) c2071123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2071123));
	wire w1991124;
	repeater #(1, 1'b1, 0, 0) c1991124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991124));
	wire w2001124;
	repeater #(1, 1'b1, 0, 0) c2001124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2001124));
	wire w1991125;
	repeater #(4, 1'b1, 0, 0) c1991125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1991125));
	wire w1861126;

	wire w1871126;

	wire w1901126;
	repeater #(1, 1'b0, 0, 0) c1901126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901126));
	wire w1911126;

	wire w1941126;

	wire w1951126;

	wire w1981126;
	repeater #(1, 1'b0, 0, 0) c1981126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1981126));
	wire w1991126;

	wire w2021126;

	wire w2031126;

	wire w2061126;
	repeater #(1, 1'b1, 0, 0) c2061126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2061126));
	wire w2071126;

	wire w2001128;
	torch #(1'b1) c2001128 (.i_clk(tick), .i_in(), .o_out(w2001128));
	wire w169046;
	repeater #(1, 1'b0, 0, 0) c169046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169046));
	wire w170047;
	repeater #(1, 1'b0, 0, 0) c170047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170047));
	wire w132048;
	repeater #(1, 1'b1, 0, 0) c132048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w132048));
	wire w149048;
	repeater #(2, 1'b1, 0, 0) c149048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w149048));
	wire w150048;
	repeater #(1, 1'b1, 0, 0) c150048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150048));
	wire w151048;

	wire w166048;

	wire w169048;
	repeater #(1, 1'b1, 0, 0) c169048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w169048));
	wire w179048;
	repeater #(1, 1'b1, 0, 0) c179048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179048));
	wire w184048;
	repeater #(1, 1'b1, 0, 0) c184048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184048));
	wire w168049;
	repeater #(1, 1'b0, 0, 0) c168049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168049));
	wire w181049;

	wire w182049;

	wire w182051;
	repeater #(1, 1'b0, 0, 0) c182051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182051));
	wire w196051;
	repeater #(1, 1'b1, 0, 0) c196051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196051));
	wire w196052;

	wire w198053;
	repeater #(1, 1'b0, 0, 0) c198053 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198053));
	wire w167054;
	repeater #(1, 1'b0, 0, 0) c167054 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167054));
	wire w130062;
	repeater #(1, 1'b1, 0, 0) c130062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130062));
	wire w198069;
	repeater #(1, 1'b0, 0, 0) c198069 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198069));
	wire w196075;
	repeater #(1, 1'b1, 0, 0) c196075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196075));
	wire w196076;

	wire w198077;
	repeater #(1, 1'b0, 0, 0) c198077 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198077));
	wire w198093;
	repeater #(1, 1'b0, 0, 0) c198093 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w198093));
	wire w196099;
	repeater #(1, 1'b1, 0, 0) c196099 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w196099));
	wire w1960100;

	wire w1980101;
	repeater #(1, 1'b0, 0, 0) c1980101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980101));
	wire w1980117;
	repeater #(1, 1'b0, 0, 0) c1980117 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980117));
	wire w1960123;
	repeater #(1, 1'b1, 0, 0) c1960123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1960123));
	wire w1960124;

	wire w1980125;
	repeater #(1, 1'b0, 0, 0) c1980125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980125));
	wire w1980141;
	repeater #(1, 1'b0, 0, 0) c1980141 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980141));
	wire w1960147;
	repeater #(1, 1'b1, 0, 0) c1960147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1960147));
	wire w1960148;

	wire w1980149;
	repeater #(1, 1'b0, 0, 0) c1980149 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980149));
	wire w1980165;
	repeater #(1, 1'b0, 0, 0) c1980165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1980165));
	wire w2000170;
	repeater #(1, 1'b0, 0, 0) c2000170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w2000170));
	wire w2010172;

	wire w2040172;
	assign outputs[123] = ();
	wire w2010173;

	wire w1990174;
	repeater #(1, 1'b0, 0, 0) c1990174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1990174));
	wire w133148;

	wire w170153;
	repeater #(1, 1'b0, 0, 0) c170153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170153));
	wire w171153;

	wire w174153;
	repeater #(1, 1'b0, 0, 0) c174153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174153));
	wire w175153;

	wire w178153;
	repeater #(1, 1'b0, 0, 0) c178153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178153));
	wire w179153;

	wire w182153;
	repeater #(1, 1'b0, 0, 0) c182153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182153));
	wire w183153;

	wire w186153;
	repeater #(1, 1'b0, 0, 0) c186153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186153));
	wire w187153;

	wire w190153;
	repeater #(1, 1'b0, 0, 0) c190153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190153));
	wire w191153;

	wire w194153;
	repeater #(1, 1'b0, 0, 0) c194153 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194153));
	wire w195153;

	wire w170156;
	repeater #(1, 1'b0, 0, 0) c170156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170156));
	wire w175156;
	repeater #(1, 1'b0, 0, 0) c175156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175156));
	wire w178156;
	repeater #(1, 1'b0, 0, 0) c178156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178156));
	wire w183156;
	repeater #(1, 1'b0, 0, 0) c183156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183156));
	wire w186156;
	repeater #(1, 1'b0, 0, 0) c186156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186156));
	wire w191156;
	repeater #(1, 1'b0, 0, 0) c191156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191156));
	wire w172157;

	wire w173157;

	wire w180157;

	wire w181157;

	wire w188157;

	wire w189157;

	wire w194157;
	repeater #(4, 1'b0, 0, 0) c194157 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194157));
	wire w170158;
	repeater #(4, 1'b0, 0, 0) c170158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170158));
	wire w175158;
	repeater #(2, 1'b0, 0, 0) c175158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175158));
	wire w178158;
	repeater #(4, 1'b0, 0, 0) c178158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178158));
	wire w183158;
	repeater #(2, 1'b0, 0, 0) c183158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183158));
	wire w186158;
	repeater #(4, 1'b0, 0, 0) c186158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186158));
	wire w191158;
	repeater #(2, 1'b0, 0, 0) c191158 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191158));
	wire w175160;
	repeater #(2, 1'b0, 0, 0) c175160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175160));
	wire w183160;
	repeater #(2, 1'b0, 0, 0) c183160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183160));
	wire w191160;
	repeater #(2, 1'b0, 0, 0) c191160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191160));
	wire w129161;

	wire w171161;
	repeater #(1, 1'b0, 0, 0) c171161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171161));
	wire w179161;
	repeater #(1, 1'b1, 0, 0) c179161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179161));
	wire w187161;
	repeater #(1, 1'b1, 0, 0) c187161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187161));
	wire w194161;
	repeater #(2, 1'b0, 0, 0) c194161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194161));
	wire w170163;

	wire w171163;

	wire w174163;
	repeater #(1, 1'b0, 0, 0) c174163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174163));
	wire w175163;

	wire w178163;

	wire w179163;

	wire w182163;
	repeater #(1, 1'b1, 0, 0) c182163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182163));
	wire w183163;

	wire w186163;

	wire w187163;

	wire w190163;
	repeater #(1, 1'b1, 0, 0) c190163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190163));
	wire w191163;

	wire w170166;
	repeater #(1, 1'b0, 0, 0) c170166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170166));
	wire w175166;
	repeater #(1, 1'b0, 0, 0) c175166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175166));
	wire w186166;
	repeater #(1, 1'b0, 0, 0) c186166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186166));
	wire w191166;
	repeater #(1, 1'b0, 0, 0) c191166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191166));
	wire w172167;

	wire w173167;

	wire w177167;
	repeater #(1, 1'b0, 0, 0) c177167 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177167));
	wire w180167;

	wire w181167;

	wire w188167;

	wire w189167;

	wire w170168;
	repeater #(4, 1'b0, 0, 0) c170168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170168));
	wire w175168;
	repeater #(2, 1'b0, 0, 0) c175168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175168));
	wire w176168;
	repeater #(1, 1'b0, 0, 0) c176168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176168));
	wire w178168;
	repeater #(4, 1'b0, 0, 0) c178168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178168));
	wire w183168;
	repeater #(1, 1'b0, 0, 0) c183168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183168));
	wire w186168;
	repeater #(4, 1'b0, 0, 0) c186168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186168));
	wire w191168;
	repeater #(2, 1'b0, 0, 0) c191168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191168));
	wire w175170;
	repeater #(2, 1'b0, 0, 0) c175170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175170));
	wire w191170;
	repeater #(2, 1'b0, 0, 0) c191170 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191170));
	wire w171171;
	repeater #(1, 1'b0, 0, 0) c171171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171171));
	wire w179171;
	repeater #(1, 1'b1, 0, 0) c179171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179171));
	wire w183171;
	repeater #(1, 1'b0, 0, 0) c183171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183171));
	wire w184171;
	repeater #(1, 1'b0, 0, 0) c184171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184171));
	wire w187171;
	repeater #(1, 1'b1, 0, 0) c187171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187171));
	wire w183172;
	repeater #(4, 1'b0, 0, 0) c183172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183172));
	wire w170173;

	wire w171173;

	wire w174173;
	repeater #(1, 1'b0, 0, 0) c174173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174173));
	wire w175173;

	wire w178173;

	wire w179173;

	wire w182173;
	repeater #(1, 1'b1, 0, 0) c182173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182173));
	wire w183173;

	wire w186173;

	wire w187173;

	wire w190173;
	repeater #(1, 1'b1, 0, 0) c190173 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190173));
	wire w191173;

	wire w184175;
	torch #(1'b0) c184175 (.i_clk(tick), .i_in(), .o_out(w184175));
	wire w170177;
	repeater #(1, 1'b1, 0, 0) c170177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170177));
	wire w171177;

	wire w174177;
	repeater #(1, 1'b1, 0, 0) c174177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174177));
	wire w175177;

	wire w178177;
	repeater #(1, 1'b1, 0, 0) c178177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178177));
	wire w179177;

	wire w182177;
	repeater #(1, 1'b1, 0, 0) c182177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182177));
	wire w183177;

	wire w186177;
	repeater #(1, 1'b1, 0, 0) c186177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186177));
	wire w187177;

	wire w190177;
	repeater #(1, 1'b1, 0, 0) c190177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190177));
	wire w191177;

	wire w194177;
	repeater #(1, 1'b1, 0, 0) c194177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194177));
	wire w195177;

	wire w170180;
	repeater #(1, 1'b1, 0, 0) c170180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170180));
	wire w175180;
	repeater #(1, 1'b1, 0, 0) c175180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175180));
	wire w178180;
	repeater #(1, 1'b1, 0, 0) c178180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178180));
	wire w183180;
	repeater #(1, 1'b1, 0, 0) c183180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183180));
	wire w186180;
	repeater #(1, 1'b1, 0, 0) c186180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186180));
	wire w191180;
	repeater #(1, 1'b1, 0, 0) c191180 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191180));
	wire w172181;

	wire w173181;

	wire w180181;

	wire w181181;

	wire w188181;

	wire w189181;

	wire w194181;
	repeater #(4, 1'b1, 0, 0) c194181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194181));
	wire w170182;
	repeater #(4, 1'b1, 0, 0) c170182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170182));
	wire w175182;
	repeater #(2, 1'b1, 0, 0) c175182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175182));
	wire w178182;
	repeater #(4, 1'b1, 0, 0) c178182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178182));
	wire w183182;
	repeater #(2, 1'b1, 0, 0) c183182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183182));
	wire w186182;
	repeater #(4, 1'b1, 0, 0) c186182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186182));
	wire w191182;
	repeater #(2, 1'b1, 0, 0) c191182 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191182));
	wire w175184;
	repeater #(2, 1'b1, 0, 0) c175184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175184));
	wire w183184;
	repeater #(2, 1'b1, 0, 0) c183184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183184));
	wire w191184;
	repeater #(2, 1'b1, 0, 0) c191184 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191184));
	wire w171185;
	repeater #(1, 1'b1, 0, 0) c171185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171185));
	wire w179185;
	repeater #(1, 1'b0, 0, 0) c179185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179185));
	wire w187185;
	repeater #(1, 1'b1, 0, 0) c187185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187185));
	wire w194185;
	repeater #(2, 1'b1, 0, 0) c194185 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w194185));
	wire w170187;

	wire w171187;

	wire w174187;
	repeater #(1, 1'b1, 0, 0) c174187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174187));
	wire w175187;

	wire w178187;

	wire w179187;

	wire w182187;
	repeater #(1, 1'b0, 0, 0) c182187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182187));
	wire w183187;

	wire w186187;

	wire w187187;

	wire w190187;
	repeater #(1, 1'b1, 0, 0) c190187 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190187));
	wire w191187;

	wire w170190;
	repeater #(1, 1'b1, 0, 0) c170190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170190));
	wire w175190;
	repeater #(1, 1'b1, 0, 0) c175190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175190));
	wire w186190;
	repeater #(1, 1'b1, 0, 0) c186190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186190));
	wire w191190;
	repeater #(1, 1'b1, 0, 0) c191190 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191190));
	wire w172191;

	wire w173191;

	wire w177191;
	repeater #(1, 1'b1, 0, 0) c177191 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w177191));
	wire w180191;

	wire w181191;

	wire w188191;

	wire w189191;

	wire w170192;
	repeater #(4, 1'b1, 0, 0) c170192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170192));
	wire w175192;
	repeater #(2, 1'b1, 0, 0) c175192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175192));
	wire w176192;
	repeater #(1, 1'b1, 0, 0) c176192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w176192));
	wire w178192;
	repeater #(4, 1'b1, 0, 0) c178192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178192));
	wire w183192;
	repeater #(1, 1'b1, 0, 0) c183192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183192));
	wire w186192;
	repeater #(4, 1'b1, 0, 0) c186192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w186192));
	wire w191192;
	repeater #(2, 1'b1, 0, 0) c191192 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191192));
	wire w175194;
	repeater #(2, 1'b1, 0, 0) c175194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175194));
	wire w191194;
	repeater #(2, 1'b1, 0, 0) c191194 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w191194));
	wire w171195;
	repeater #(1, 1'b0, 0, 0) c171195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171195));
	wire w179195;
	repeater #(1, 1'b1, 0, 0) c179195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w179195));
	wire w183195;
	repeater #(1, 1'b1, 0, 0) c183195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183195));
	wire w184195;
	repeater #(1, 1'b1, 0, 0) c184195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184195));
	wire w187195;
	repeater #(1, 1'b1, 0, 0) c187195 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w187195));
	wire w183196;
	repeater #(4, 1'b1, 0, 0) c183196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183196));
	wire w170197;

	wire w171197;

	wire w174197;
	repeater #(1, 1'b0, 0, 0) c174197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174197));
	wire w175197;

	wire w178197;

	wire w179197;

	wire w182197;
	repeater #(1, 1'b1, 0, 0) c182197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182197));
	wire w183197;

	wire w186197;

	wire w187197;

	wire w190197;
	repeater #(1, 1'b1, 0, 0) c190197 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w190197));
	wire w191197;

	wire w184199;
	torch #(1'b1) c184199 (.i_clk(tick), .i_in(), .o_out(w184199));
	wire w1701101;
	repeater #(1, 1'b0, 0, 0) c1701101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701101));
	wire w1711101;

	wire w1741101;
	repeater #(1, 1'b0, 0, 0) c1741101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741101));
	wire w1751101;

	wire w1781101;
	repeater #(1, 1'b0, 0, 0) c1781101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781101));
	wire w1791101;

	wire w1821101;
	repeater #(1, 1'b0, 0, 0) c1821101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821101));
	wire w1831101;

	wire w1861101;
	repeater #(1, 1'b0, 0, 0) c1861101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861101));
	wire w1871101;

	wire w1901101;
	repeater #(1, 1'b1, 0, 0) c1901101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901101));
	wire w1911101;

	wire w1941101;
	repeater #(1, 1'b1, 0, 0) c1941101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941101));
	wire w1951101;

	wire w1701104;
	repeater #(1, 1'b0, 0, 0) c1701104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701104));
	wire w1751104;
	repeater #(1, 1'b0, 0, 0) c1751104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751104));
	wire w1781104;
	repeater #(1, 1'b0, 0, 0) c1781104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781104));
	wire w1831104;
	repeater #(1, 1'b0, 0, 0) c1831104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831104));
	wire w1861104;
	repeater #(1, 1'b0, 0, 0) c1861104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861104));
	wire w1911104;
	repeater #(1, 1'b1, 0, 0) c1911104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911104));
	wire w1721105;

	wire w1731105;

	wire w1801105;

	wire w1811105;

	wire w1881105;

	wire w1891105;

	wire w1941105;
	repeater #(4, 1'b1, 0, 0) c1941105 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941105));
	wire w1701106;
	repeater #(4, 1'b0, 0, 0) c1701106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701106));
	wire w1751106;
	repeater #(2, 1'b0, 0, 0) c1751106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751106));
	wire w1781106;
	repeater #(4, 1'b0, 0, 0) c1781106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781106));
	wire w1831106;
	repeater #(2, 1'b0, 0, 0) c1831106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831106));
	wire w1861106;
	repeater #(4, 1'b0, 0, 0) c1861106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861106));
	wire w1911106;
	repeater #(2, 1'b1, 0, 0) c1911106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911106));
	wire w1751108;
	repeater #(2, 1'b0, 0, 0) c1751108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751108));
	wire w1831108;
	repeater #(2, 1'b0, 0, 0) c1831108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831108));
	wire w1911108;
	repeater #(2, 1'b1, 0, 0) c1911108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911108));
	wire w1711109;
	repeater #(1, 1'b0, 0, 0) c1711109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1711109));
	wire w1791109;
	repeater #(1, 1'b0, 0, 0) c1791109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1791109));
	wire w1871109;
	repeater #(1, 1'b1, 0, 0) c1871109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1871109));
	wire w1941109;
	repeater #(2, 1'b1, 0, 0) c1941109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941109));
	wire w1701111;

	wire w1711111;

	wire w1741111;
	repeater #(1, 1'b0, 0, 0) c1741111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741111));
	wire w1751111;

	wire w1781111;

	wire w1791111;

	wire w1821111;
	repeater #(1, 1'b0, 0, 0) c1821111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821111));
	wire w1831111;

	wire w1861111;

	wire w1871111;

	wire w1901111;
	repeater #(1, 1'b1, 0, 0) c1901111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901111));
	wire w1911111;

	wire w1701114;
	repeater #(1, 1'b0, 0, 0) c1701114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701114));
	wire w1751114;
	repeater #(1, 1'b0, 0, 0) c1751114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751114));
	wire w1861114;
	repeater #(1, 1'b0, 0, 0) c1861114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861114));
	wire w1911114;
	repeater #(1, 1'b1, 0, 0) c1911114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911114));
	wire w1721115;

	wire w1731115;

	wire w1771115;
	repeater #(1, 1'b0, 0, 0) c1771115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1771115));
	wire w1801115;

	wire w1811115;

	wire w1881115;

	wire w1891115;

	wire w1701116;
	repeater #(4, 1'b0, 0, 0) c1701116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701116));
	wire w1751116;
	repeater #(2, 1'b0, 0, 0) c1751116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751116));
	wire w1761116;
	repeater #(1, 1'b0, 0, 0) c1761116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1761116));
	wire w1781116;
	repeater #(4, 1'b0, 0, 0) c1781116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781116));
	wire w1831116;
	repeater #(1, 1'b0, 0, 0) c1831116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831116));
	wire w1861116;
	repeater #(4, 1'b0, 0, 0) c1861116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861116));
	wire w1911116;
	repeater #(2, 1'b1, 0, 0) c1911116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911116));
	wire w1751118;
	repeater #(2, 1'b0, 0, 0) c1751118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751118));
	wire w1911118;
	repeater #(2, 1'b1, 0, 0) c1911118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911118));
	wire w1711119;
	repeater #(1, 1'b0, 0, 0) c1711119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1711119));
	wire w1791119;
	repeater #(1, 1'b1, 0, 0) c1791119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1791119));
	wire w1831119;
	repeater #(1, 1'b0, 0, 0) c1831119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831119));
	wire w1841119;
	repeater #(1, 1'b0, 0, 0) c1841119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1841119));
	wire w1871119;
	repeater #(1, 1'b1, 0, 0) c1871119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1871119));
	wire w1831120;
	repeater #(4, 1'b0, 0, 0) c1831120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831120));
	wire w1701121;

	wire w1711121;

	wire w1741121;
	repeater #(1, 1'b0, 0, 0) c1741121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741121));
	wire w1751121;

	wire w1781121;

	wire w1791121;

	wire w1821121;
	repeater #(1, 1'b1, 0, 0) c1821121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821121));
	wire w1831121;

	wire w1861121;

	wire w1871121;

	wire w1901121;
	repeater #(1, 1'b1, 0, 0) c1901121 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901121));
	wire w1911121;

	wire w1841123;
	torch #(1'b0) c1841123 (.i_clk(tick), .i_in(), .o_out(w1841123));
	wire w1701125;
	repeater #(1, 1'b0, 0, 0) c1701125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701125));
	wire w1711125;

	wire w1741125;
	repeater #(1, 1'b0, 0, 0) c1741125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741125));
	wire w1751125;

	wire w1781125;
	repeater #(1, 1'b0, 0, 0) c1781125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781125));
	wire w1791125;

	wire w1821125;
	repeater #(1, 1'b0, 0, 0) c1821125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821125));
	wire w1831125;

	wire w1861125;
	repeater #(1, 1'b0, 0, 0) c1861125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861125));
	wire w1871125;

	wire w1901125;
	repeater #(1, 1'b0, 0, 0) c1901125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901125));
	wire w1911125;

	wire w1941125;
	repeater #(1, 1'b0, 0, 0) c1941125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941125));
	wire w1951125;

	wire w1701128;
	repeater #(1, 1'b0, 0, 0) c1701128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701128));
	wire w1751128;
	repeater #(1, 1'b0, 0, 0) c1751128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751128));
	wire w1781128;
	repeater #(1, 1'b0, 0, 0) c1781128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781128));
	wire w1831128;
	repeater #(1, 1'b0, 0, 0) c1831128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831128));
	wire w1861128;
	repeater #(1, 1'b0, 0, 0) c1861128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861128));
	wire w1911128;
	repeater #(1, 1'b0, 0, 0) c1911128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911128));
	wire w1721129;

	wire w1731129;

	wire w1801129;

	wire w1811129;

	wire w1881129;

	wire w1891129;

	wire w1941129;
	repeater #(4, 1'b0, 0, 0) c1941129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941129));
	wire w1701130;
	repeater #(4, 1'b0, 0, 0) c1701130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701130));
	wire w1751130;
	repeater #(2, 1'b0, 0, 0) c1751130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751130));
	wire w1781130;
	repeater #(4, 1'b0, 0, 0) c1781130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781130));
	wire w1831130;
	repeater #(2, 1'b0, 0, 0) c1831130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831130));
	wire w1861130;
	repeater #(4, 1'b0, 0, 0) c1861130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1861130));
	wire w1911130;
	repeater #(2, 1'b0, 0, 0) c1911130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911130));
	wire w1751132;
	repeater #(2, 1'b0, 0, 0) c1751132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751132));
	wire w1831132;
	repeater #(2, 1'b0, 0, 0) c1831132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1831132));
	wire w1911132;
	repeater #(2, 1'b0, 0, 0) c1911132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1911132));
	wire w1711133;
	repeater #(1, 1'b0, 0, 0) c1711133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1711133));
	wire w1791133;
	repeater #(1, 1'b0, 0, 0) c1791133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1791133));
	wire w1871133;
	repeater #(1, 1'b0, 0, 0) c1871133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1871133));
	wire w1941133;
	repeater #(2, 1'b0, 0, 0) c1941133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1941133));
	wire w1701135;

	wire w1711135;

	wire w1741135;
	repeater #(1, 1'b0, 0, 0) c1741135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741135));
	wire w1751135;

	wire w1781135;

	wire w1791135;

	wire w1821135;
	repeater #(1, 1'b0, 0, 0) c1821135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1821135));
	wire w1831135;

	wire w1861135;

	wire w1871135;

	wire w1901135;
	repeater #(1, 1'b0, 0, 0) c1901135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1901135));
	wire w1911135;

	wire w15402;
	repeater #(1, 1'b0, 0, 0) c15402 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15402));
	wire w15902;
	repeater #(1, 1'b0, 0, 0) c15902 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15902));
	wire w17002;
	repeater #(1, 1'b0, 0, 0) c17002 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17002));
	wire w17502;
	repeater #(1, 1'b0, 0, 0) c17502 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17502));
	wire w15603;

	wire w15703;

	wire w16103;
	repeater #(1, 1'b0, 0, 0) c16103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16103));
	wire w16403;

	wire w16503;

	wire w17203;

	wire w17303;

	wire w15404;
	repeater #(4, 1'b0, 0, 0) c15404 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15404));
	wire w15904;
	repeater #(2, 1'b0, 0, 0) c15904 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15904));
	wire w16004;
	repeater #(1, 1'b0, 0, 0) c16004 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16004));
	wire w16204;
	repeater #(4, 1'b0, 0, 0) c16204 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16204));
	wire w16704;
	repeater #(1, 1'b0, 0, 0) c16704 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16704));
	wire w17004;
	repeater #(4, 1'b0, 0, 0) c17004 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17004));
	wire w17504;
	repeater #(2, 1'b0, 0, 0) c17504 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17504));
	wire w15906;
	repeater #(2, 1'b0, 0, 0) c15906 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15906));
	wire w17506;
	repeater #(2, 1'b0, 0, 0) c17506 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17506));
	wire w15507;
	repeater #(1, 1'b0, 0, 0) c15507 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15507));
	wire w16307;
	repeater #(1, 1'b0, 0, 0) c16307 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16307));
	wire w16707;
	repeater #(1, 1'b0, 0, 0) c16707 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16707));
	wire w16807;
	repeater #(1, 1'b0, 0, 0) c16807 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16807));
	wire w17107;
	repeater #(1, 1'b0, 0, 0) c17107 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17107));
	wire w16708;
	repeater #(4, 1'b0, 0, 0) c16708 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16708));
	wire w15409;

	wire w15509;

	wire w15809;
	repeater #(1, 1'b0, 0, 0) c15809 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15809));
	wire w15909;

	wire w16209;

	wire w16309;

	wire w16609;
	repeater #(1, 1'b0, 0, 0) c16609 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16609));
	wire w16709;

	wire w17009;

	wire w17109;

	wire w17409;
	repeater #(1, 1'b0, 0, 0) c17409 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17409));
	wire w17509;

	wire w168011;
	torch #(1'b0) c168011 (.i_clk(tick), .i_in(), .o_out(w168011));
	wire w154013;
	repeater #(1, 1'b1, 0, 0) c154013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154013));
	wire w155013;

	wire w158013;
	repeater #(1, 1'b1, 0, 0) c158013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158013));
	wire w159013;

	wire w162013;
	repeater #(1, 1'b1, 0, 0) c162013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162013));
	wire w163013;

	wire w166013;
	repeater #(1, 1'b1, 0, 0) c166013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166013));
	wire w167013;

	wire w170013;
	repeater #(1, 1'b1, 0, 0) c170013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170013));
	wire w171013;

	wire w174013;
	repeater #(1, 1'b1, 0, 0) c174013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174013));
	wire w175013;

	wire w178013;
	repeater #(1, 1'b0, 0, 0) c178013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178013));
	wire w179013;

	wire w154016;
	repeater #(1, 1'b1, 0, 0) c154016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154016));
	wire w159016;
	repeater #(1, 1'b1, 0, 0) c159016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159016));
	wire w162016;
	repeater #(1, 1'b1, 0, 0) c162016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162016));
	wire w167016;
	repeater #(1, 1'b1, 0, 0) c167016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167016));
	wire w170016;
	repeater #(1, 1'b1, 0, 0) c170016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170016));
	wire w175016;
	repeater #(1, 1'b1, 0, 0) c175016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175016));
	wire w156017;

	wire w157017;

	wire w164017;

	wire w165017;

	wire w172017;

	wire w173017;

	wire w178017;
	repeater #(4, 1'b0, 0, 0) c178017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178017));
	wire w154018;
	repeater #(4, 1'b1, 0, 0) c154018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154018));
	wire w159018;
	repeater #(2, 1'b1, 0, 0) c159018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159018));
	wire w162018;
	repeater #(4, 1'b1, 0, 0) c162018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162018));
	wire w167018;
	repeater #(2, 1'b1, 0, 0) c167018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167018));
	wire w170018;
	repeater #(4, 1'b1, 0, 0) c170018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170018));
	wire w175018;
	repeater #(2, 1'b1, 0, 0) c175018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175018));
	wire w159020;
	repeater #(2, 1'b1, 0, 0) c159020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159020));
	wire w167020;
	repeater #(2, 1'b1, 0, 0) c167020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167020));
	wire w175020;
	repeater #(2, 1'b1, 0, 0) c175020 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175020));
	wire w155021;
	repeater #(1, 1'b0, 0, 0) c155021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155021));
	wire w163021;
	repeater #(1, 1'b0, 0, 0) c163021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163021));
	wire w171021;
	repeater #(1, 1'b0, 0, 0) c171021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171021));
	wire w178021;
	repeater #(2, 1'b0, 0, 0) c178021 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178021));
	wire w154023;

	wire w155023;

	wire w158023;
	repeater #(1, 1'b0, 0, 0) c158023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158023));
	wire w159023;

	wire w162023;

	wire w163023;

	wire w166023;
	repeater #(1, 1'b0, 0, 0) c166023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166023));
	wire w167023;

	wire w170023;

	wire w171023;

	wire w174023;
	repeater #(1, 1'b0, 0, 0) c174023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174023));
	wire w175023;

	wire w154026;
	repeater #(1, 1'b1, 0, 0) c154026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154026));
	wire w159026;
	repeater #(1, 1'b1, 0, 0) c159026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159026));
	wire w170026;
	repeater #(1, 1'b1, 0, 0) c170026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170026));
	wire w175026;
	repeater #(1, 1'b0, 0, 0) c175026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175026));
	wire w156027;

	wire w157027;

	wire w161027;
	repeater #(1, 1'b1, 0, 0) c161027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w161027));
	wire w164027;

	wire w165027;

	wire w172027;

	wire w173027;

	wire w154028;
	repeater #(4, 1'b1, 0, 0) c154028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154028));
	wire w159028;
	repeater #(2, 1'b1, 0, 0) c159028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159028));
	wire w160028;
	repeater #(1, 1'b1, 0, 0) c160028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w160028));
	wire w162028;
	repeater #(4, 1'b1, 0, 0) c162028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162028));
	wire w167028;
	repeater #(1, 1'b1, 0, 0) c167028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167028));
	wire w170028;
	repeater #(4, 1'b1, 0, 0) c170028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170028));
	wire w175028;
	repeater #(2, 1'b0, 0, 0) c175028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175028));
	wire w159030;
	repeater #(2, 1'b1, 0, 0) c159030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159030));
	wire w175030;
	repeater #(2, 1'b0, 0, 0) c175030 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w175030));
	wire w155031;
	repeater #(1, 1'b0, 0, 0) c155031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155031));
	wire w163031;
	repeater #(1, 1'b0, 0, 0) c163031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163031));
	wire w167031;
	repeater #(1, 1'b1, 0, 0) c167031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167031));
	wire w168031;
	repeater #(1, 1'b1, 0, 0) c168031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168031));
	wire w171031;
	repeater #(1, 1'b1, 0, 0) c171031 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171031));
	wire w167032;
	repeater #(4, 1'b1, 0, 0) c167032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167032));
	wire w154033;

	wire w155033;

	wire w158033;
	repeater #(1, 1'b0, 0, 0) c158033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158033));
	wire w159033;

	wire w162033;

	wire w163033;

	wire w166033;
	repeater #(1, 1'b0, 0, 0) c166033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166033));
	wire w167033;

	wire w170033;

	wire w171033;

	wire w174033;
	repeater #(1, 1'b1, 0, 0) c174033 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174033));
	wire w175033;

	wire w168035;
	torch #(1'b1) c168035 (.i_clk(tick), .i_in(), .o_out(w168035));
	wire w153089;
	repeater #(1, 1'b0, 0, 0) c153089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153089));
	wire w154090;
	repeater #(1, 1'b0, 0, 0) c154090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154090));
	wire w116091;
	repeater #(1, 1'b1, 0, 0) c116091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w116091));
	wire w133091;
	repeater #(2, 1'b1, 0, 0) c133091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w133091));
	wire w134091;
	repeater #(1, 1'b1, 0, 0) c134091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134091));
	wire w135091;

	wire w150091;

	wire w153091;
	repeater #(1, 1'b1, 0, 0) c153091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w153091));
	wire w163091;
	repeater #(1, 1'b1, 0, 0) c163091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163091));
	wire w168091;
	repeater #(1, 1'b1, 0, 0) c168091 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168091));
	wire w152092;
	repeater #(1, 1'b0, 0, 0) c152092 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152092));
	wire w165092;

	wire w166092;

	wire w166094;
	repeater #(1, 1'b0, 0, 0) c166094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166094));
	wire w180094;
	repeater #(1, 1'b1, 0, 0) c180094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180094));
	wire w180095;

	wire w182096;
	repeater #(1, 1'b0, 0, 0) c182096 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182096));
	wire w151097;
	repeater #(1, 1'b0, 0, 0) c151097 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151097));
	wire w1550102;
	repeater #(1, 1'b0, 0, 0) c1550102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550102));
	wire w1630102;
	repeater #(1, 1'b0, 0, 0) c1630102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630102));
	wire w1710102;
	repeater #(1, 1'b0, 0, 0) c1710102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710102));
	wire w1560103;

	wire w1640103;

	wire w1720103;

	wire w1550112;
	repeater #(1, 1'b0, 0, 0) c1550112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550112));
	wire w1630112;
	repeater #(1, 1'b0, 0, 0) c1630112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630112));
	wire w1710112;
	repeater #(1, 1'b0, 0, 0) c1710112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710112));
	wire w1820112;
	repeater #(1, 1'b0, 0, 0) c1820112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820112));
	wire w1560113;

	wire w1640113;

	wire w1720113;

	wire w1800118;
	repeater #(1, 1'b1, 0, 0) c1800118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800118));
	wire w1800119;

	wire w1820120;
	repeater #(1, 1'b0, 0, 0) c1820120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820120));
	wire w1550126;
	repeater #(1, 1'b0, 0, 0) c1550126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550126));
	wire w1630126;
	repeater #(1, 1'b0, 0, 0) c1630126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630126));
	wire w1710126;
	repeater #(1, 1'b0, 0, 0) c1710126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710126));
	wire w1560127;

	wire w1640127;

	wire w1720127;

	wire w1550136;
	repeater #(1, 1'b0, 0, 0) c1550136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550136));
	wire w1630136;
	repeater #(1, 1'b0, 0, 0) c1630136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630136));
	wire w1710136;
	repeater #(1, 1'b0, 0, 0) c1710136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710136));
	wire w1820136;
	repeater #(1, 1'b0, 0, 0) c1820136 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820136));
	wire w1560137;

	wire w1640137;

	wire w1720137;

	wire w1800142;
	repeater #(1, 1'b1, 0, 0) c1800142 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800142));
	wire w1800143;

	wire w1820144;
	repeater #(1, 1'b0, 0, 0) c1820144 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820144));
	wire w1550150;
	repeater #(1, 1'b0, 0, 0) c1550150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550150));
	wire w1630150;
	repeater #(1, 1'b0, 0, 0) c1630150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630150));
	wire w1710150;
	repeater #(1, 1'b0, 0, 0) c1710150 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710150));
	wire w1560151;

	wire w1640151;

	wire w1720151;

	wire w1550160;
	repeater #(1, 1'b0, 0, 0) c1550160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550160));
	wire w1630160;
	repeater #(1, 1'b0, 0, 0) c1630160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630160));
	wire w1710160;
	repeater #(1, 1'b0, 0, 0) c1710160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710160));
	wire w1820160;
	repeater #(1, 1'b0, 0, 0) c1820160 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820160));
	wire w1560161;

	wire w1640161;

	wire w1720161;

	wire w1800166;
	repeater #(1, 1'b1, 0, 0) c1800166 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1800166));
	wire w1800167;

	wire w1820168;
	repeater #(1, 1'b0, 0, 0) c1820168 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1820168));
	wire w1550174;
	repeater #(1, 1'b0, 0, 0) c1550174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550174));
	wire w1630174;
	repeater #(1, 1'b0, 0, 0) c1630174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1630174));
	wire w1710174;
	repeater #(1, 1'b0, 0, 0) c1710174 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1710174));
	wire w1560175;

	wire w1640175;

	wire w1720175;

	wire w15515;
	repeater #(1, 1'b0, 0, 0) c15515 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15515));
	wire w16315;
	repeater #(1, 1'b0, 0, 0) c16315 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16315));
	wire w17115;
	repeater #(1, 1'b0, 0, 0) c17115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w17115));
	wire w18215;
	repeater #(1, 1'b0, 0, 0) c18215 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w18215));
	wire w15616;

	wire w16416;

	wire w17216;

	wire w180111;
	repeater #(1, 1'b1, 0, 0) c180111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w180111));
	wire w180112;

	wire w182113;
	repeater #(1, 1'b0, 0, 0) c182113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182113));
	wire w155119;
	repeater #(1, 1'b0, 0, 0) c155119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155119));
	wire w163119;
	repeater #(1, 1'b0, 0, 0) c163119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163119));
	wire w171119;
	repeater #(1, 1'b0, 0, 0) c171119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171119));
	wire w156120;

	wire w164120;

	wire w172120;

	wire w155129;
	repeater #(1, 1'b0, 0, 0) c155129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155129));
	wire w163129;
	repeater #(1, 1'b0, 0, 0) c163129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w163129));
	wire w171129;
	repeater #(1, 1'b0, 0, 0) c171129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w171129));
	wire w182129;
	repeater #(1, 1'b0, 0, 0) c182129 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w182129));
	wire w156130;

	wire w164130;

	wire w172130;

	wire w184134;
	repeater #(1, 1'b0, 0, 0) c184134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w184134));
	wire w185136;

	wire w188136;
	assign outputs[124] = ();
	wire w185137;

	wire w183138;
	repeater #(1, 1'b0, 0, 0) c183138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w183138));
	wire w154140;
	repeater #(1, 1'b0, 0, 0) c154140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154140));
	wire w158140;
	repeater #(1, 1'b0, 0, 0) c158140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158140));
	wire w162140;
	repeater #(1, 1'b0, 0, 0) c162140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162140));
	wire w166140;
	repeater #(1, 1'b0, 0, 0) c166140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166140));
	wire w170140;
	repeater #(1, 1'b0, 0, 0) c170140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170140));
	wire w174140;
	repeater #(1, 1'b0, 0, 0) c174140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174140));
	wire w178140;
	repeater #(1, 1'b0, 0, 0) c178140 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178140));
	wire w117191;

	wire w154196;
	repeater #(1, 1'b0, 0, 0) c154196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154196));
	wire w155196;

	wire w158196;
	repeater #(1, 1'b0, 0, 0) c158196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158196));
	wire w159196;

	wire w162196;
	repeater #(1, 1'b0, 0, 0) c162196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162196));
	wire w163196;

	wire w166196;
	repeater #(1, 1'b0, 0, 0) c166196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166196));
	wire w167196;

	wire w170196;
	repeater #(1, 1'b0, 0, 0) c170196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w170196));
	wire w171196;

	wire w174196;
	repeater #(1, 1'b0, 0, 0) c174196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w174196));
	wire w175196;

	wire w178196;
	repeater #(1, 1'b0, 0, 0) c178196 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w178196));
	wire w179196;

	wire w1541100;
	repeater #(1, 1'b0, 0, 0) c1541100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541100));
	wire w1621100;
	repeater #(1, 1'b0, 0, 0) c1621100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621100));
	wire w1701100;
	repeater #(1, 1'b0, 0, 0) c1701100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701100));
	wire w1781100;
	repeater #(4, 1'b0, 0, 0) c1781100 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781100));
	wire w1541101;
	repeater #(4, 1'b0, 0, 0) c1541101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541101));
	wire w1561101;

	wire w1571101;

	wire w1591101;
	repeater #(2, 1'b0, 0, 0) c1591101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591101));
	wire w1621101;
	repeater #(4, 1'b0, 0, 0) c1621101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621101));
	wire w1641101;

	wire w1651101;

	wire w1671101;
	repeater #(2, 1'b0, 0, 0) c1671101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671101));
	wire w1701101;
	repeater #(4, 1'b0, 0, 0) c1701101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701101));
	wire w1721101;

	wire w1731101;

	wire w1751101;
	repeater #(2, 1'b0, 0, 0) c1751101 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751101));
	wire w1591102;
	repeater #(1, 1'b0, 0, 0) c1591102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591102));
	wire w1671102;
	repeater #(1, 1'b0, 0, 0) c1671102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671102));
	wire w1751102;
	repeater #(1, 1'b0, 0, 0) c1751102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751102));
	wire w1591103;
	repeater #(2, 1'b0, 0, 0) c1591103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591103));
	wire w1671103;
	repeater #(2, 1'b0, 0, 0) c1671103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671103));
	wire w1751103;
	repeater #(2, 1'b0, 0, 0) c1751103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751103));
	wire w1781104;
	repeater #(2, 1'b0, 0, 0) c1781104 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781104));
	wire w1541106;

	wire w1551106;

	wire w1581106;
	repeater #(1, 1'b0, 0, 0) c1581106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581106));
	wire w1591106;

	wire w1621106;

	wire w1631106;

	wire w1661106;
	repeater #(1, 1'b1, 0, 0) c1661106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661106));
	wire w1671106;

	wire w1701106;

	wire w1711106;

	wire w1741106;
	repeater #(1, 1'b1, 0, 0) c1741106 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741106));
	wire w1751106;

	wire w1541110;
	repeater #(1, 1'b0, 0, 0) c1541110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541110));
	wire w1591110;
	repeater #(1, 1'b0, 0, 0) c1591110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591110));
	wire w1701110;
	repeater #(1, 1'b0, 0, 0) c1701110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701110));
	wire w1561111;

	wire w1571111;

	wire w1601111;
	repeater #(1, 1'b0, 0, 0) c1601111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1601111));
	wire w1621111;
	repeater #(4, 1'b0, 0, 0) c1621111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621111));
	wire w1641111;

	wire w1651111;

	wire w1701111;
	repeater #(4, 1'b0, 0, 0) c1701111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701111));
	wire w1721111;

	wire w1731111;

	wire w1751111;
	repeater #(2, 1'b0, 0, 0) c1751111 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751111));
	wire w1621112;
	repeater #(1, 1'b0, 0, 0) c1621112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621112));
	wire w1751112;
	repeater #(1, 1'b0, 0, 0) c1751112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751112));
	wire w1591113;
	repeater #(2, 1'b0, 0, 0) c1591113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591113));
	wire w1751113;
	repeater #(2, 1'b0, 0, 0) c1751113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751113));
	wire w1591114;
	repeater #(3, 1'b0, 0, 0) c1591114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591114));
	wire w1671114;
	repeater #(1, 1'b0, 0, 0) c1671114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671114));
	wire w1681114;
	repeater #(1, 1'b0, 0, 0) c1681114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1681114));
	wire w1671115;
	repeater #(4, 1'b0, 0, 0) c1671115 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671115));
	wire w1541116;

	wire w1551116;

	wire w1581116;
	repeater #(1, 1'b0, 0, 0) c1581116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581116));
	wire w1591116;

	wire w1621116;

	wire w1631116;

	wire w1661116;
	repeater #(1, 1'b1, 0, 0) c1661116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661116));
	wire w1671116;

	wire w1701116;

	wire w1711116;

	wire w1741116;
	repeater #(1, 1'b1, 0, 0) c1741116 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741116));
	wire w1751116;

	wire w1681118;
	torch #(1'b0) c1681118 (.i_clk(tick), .i_in(), .o_out(w1681118));
	wire w1541120;
	repeater #(1, 1'b1, 0, 0) c1541120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541120));
	wire w1551120;

	wire w1581120;
	repeater #(1, 1'b1, 0, 0) c1581120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581120));
	wire w1591120;

	wire w1621120;
	repeater #(1, 1'b1, 0, 0) c1621120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621120));
	wire w1631120;

	wire w1661120;
	repeater #(1, 1'b1, 0, 0) c1661120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661120));
	wire w1671120;

	wire w1701120;
	repeater #(1, 1'b1, 0, 0) c1701120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701120));
	wire w1711120;

	wire w1741120;
	repeater #(1, 1'b1, 0, 0) c1741120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741120));
	wire w1751120;

	wire w1781120;
	repeater #(1, 1'b1, 0, 0) c1781120 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781120));
	wire w1791120;

	wire w1541124;
	repeater #(1, 1'b1, 0, 0) c1541124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541124));
	wire w1621124;
	repeater #(1, 1'b1, 0, 0) c1621124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621124));
	wire w1701124;
	repeater #(1, 1'b1, 0, 0) c1701124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701124));
	wire w1781124;
	repeater #(4, 1'b1, 0, 0) c1781124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781124));
	wire w1541125;
	repeater #(4, 1'b1, 0, 0) c1541125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541125));
	wire w1561125;

	wire w1571125;

	wire w1591125;
	repeater #(2, 1'b1, 0, 0) c1591125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591125));
	wire w1621125;
	repeater #(4, 1'b1, 0, 0) c1621125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621125));
	wire w1641125;

	wire w1651125;

	wire w1671125;
	repeater #(2, 1'b1, 0, 0) c1671125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671125));
	wire w1701125;
	repeater #(4, 1'b1, 0, 0) c1701125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701125));
	wire w1721125;

	wire w1731125;

	wire w1751125;
	repeater #(2, 1'b1, 0, 0) c1751125 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751125));
	wire w1591126;
	repeater #(1, 1'b1, 0, 0) c1591126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591126));
	wire w1671126;
	repeater #(1, 1'b1, 0, 0) c1671126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671126));
	wire w1751126;
	repeater #(1, 1'b1, 0, 0) c1751126 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751126));
	wire w1591127;
	repeater #(2, 1'b1, 0, 0) c1591127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591127));
	wire w1671127;
	repeater #(2, 1'b1, 0, 0) c1671127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1671127));
	wire w1751127;
	repeater #(2, 1'b1, 0, 0) c1751127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751127));
	wire w1781128;
	repeater #(2, 1'b1, 0, 0) c1781128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1781128));
	wire w1541130;

	wire w1551130;

	wire w1581130;
	repeater #(1, 1'b1, 0, 0) c1581130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1581130));
	wire w1591130;

	wire w1621130;

	wire w1631130;

	wire w1661130;
	repeater #(1, 1'b0, 0, 0) c1661130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1661130));
	wire w1671130;

	wire w1701130;

	wire w1711130;

	wire w1741130;
	repeater #(1, 1'b1, 0, 0) c1741130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1741130));
	wire w1751130;

	wire w1541134;
	repeater #(1, 1'b1, 0, 0) c1541134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1541134));
	wire w1591134;
	repeater #(1, 1'b1, 0, 0) c1591134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1591134));
	wire w1701134;
	repeater #(1, 1'b1, 0, 0) c1701134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701134));
	wire w1561135;

	wire w1571135;

	wire w1601135;
	repeater #(1, 1'b1, 0, 0) c1601135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1601135));
	wire w1621135;
	repeater #(4, 1'b1, 0, 0) c1621135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1621135));
	wire w1641135;

	wire w1651135;

	wire w1701135;
	repeater #(4, 1'b1, 0, 0) c1701135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1701135));
	wire w1721135;

	wire w1731135;

	wire w1751135;
	repeater #(2, 1'b1, 0, 0) c1751135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1751135));
	wire w14600;
	repeater #(1, 1'b1, 0, 0) c14600 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14600));
	wire w15900;
	repeater #(1, 1'b1, 0, 0) c15900 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15900));
	wire w14301;
	repeater #(2, 1'b1, 0, 0) c14301 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14301));
	wire w15901;
	repeater #(2, 1'b1, 0, 0) c15901 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15901));
	wire w14302;
	repeater #(3, 1'b1, 0, 0) c14302 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14302));
	wire w15102;
	repeater #(1, 1'b1, 0, 0) c15102 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15102));
	wire w15202;
	repeater #(1, 1'b1, 0, 0) c15202 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15202));
	wire w15103;
	repeater #(4, 1'b1, 0, 0) c15103 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15103));
	wire w13804;

	wire w13904;

	wire w14204;
	repeater #(1, 1'b0, 0, 0) c14204 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14204));
	wire w14304;

	wire w14604;

	wire w14704;

	wire w15004;
	repeater #(1, 1'b1, 0, 0) c15004 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15004));
	wire w15104;

	wire w15404;

	wire w15504;

	wire w15804;
	repeater #(1, 1'b1, 0, 0) c15804 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15804));
	wire w15904;

	wire w15206;
	torch #(1'b1) c15206 (.i_clk(tick), .i_in(), .o_out(w15206));
	wire w13808;
	repeater #(1, 1'b0, 0, 0) c13808 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w13808));
	wire w13908;

	wire w14208;
	repeater #(1, 1'b0, 0, 0) c14208 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14208));
	wire w14308;

	wire w14608;
	repeater #(1, 1'b0, 0, 0) c14608 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14608));
	wire w14708;

	wire w15008;
	repeater #(1, 1'b0, 0, 0) c15008 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15008));
	wire w15108;

	wire w15408;
	repeater #(1, 1'b0, 0, 0) c15408 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15408));
	wire w15508;

	wire w15808;
	repeater #(1, 1'b1, 0, 0) c15808 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15808));
	wire w15908;

	wire w16208;
	repeater #(1, 1'b1, 0, 0) c16208 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16208));
	wire w16308;

	wire w138012;
	repeater #(1, 1'b0, 0, 0) c138012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138012));
	wire w146012;
	repeater #(1, 1'b0, 0, 0) c146012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146012));
	wire w154012;
	repeater #(1, 1'b0, 0, 0) c154012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154012));
	wire w162012;
	repeater #(4, 1'b1, 0, 0) c162012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162012));
	wire w138013;
	repeater #(4, 1'b0, 0, 0) c138013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138013));
	wire w140013;

	wire w141013;

	wire w143013;
	repeater #(2, 1'b0, 0, 0) c143013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143013));
	wire w146013;
	repeater #(4, 1'b0, 0, 0) c146013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146013));
	wire w148013;

	wire w149013;

	wire w151013;
	repeater #(2, 1'b0, 0, 0) c151013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151013));
	wire w154013;
	repeater #(4, 1'b0, 0, 0) c154013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154013));
	wire w156013;

	wire w157013;

	wire w159013;
	repeater #(2, 1'b1, 0, 0) c159013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159013));
	wire w143014;
	repeater #(1, 1'b0, 0, 0) c143014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143014));
	wire w151014;
	repeater #(1, 1'b0, 0, 0) c151014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151014));
	wire w159014;
	repeater #(1, 1'b1, 0, 0) c159014 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159014));
	wire w143015;
	repeater #(2, 1'b0, 0, 0) c143015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143015));
	wire w151015;
	repeater #(2, 1'b0, 0, 0) c151015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151015));
	wire w159015;
	repeater #(2, 1'b1, 0, 0) c159015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159015));
	wire w162016;
	repeater #(2, 1'b1, 0, 0) c162016 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162016));
	wire w138018;

	wire w139018;

	wire w142018;
	repeater #(1, 1'b0, 0, 0) c142018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142018));
	wire w143018;

	wire w146018;

	wire w147018;

	wire w150018;
	repeater #(1, 1'b0, 0, 0) c150018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150018));
	wire w151018;

	wire w154018;

	wire w155018;

	wire w158018;
	repeater #(1, 1'b1, 0, 0) c158018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158018));
	wire w159018;

	wire w138022;
	repeater #(1, 1'b0, 0, 0) c138022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138022));
	wire w143022;
	repeater #(1, 1'b0, 0, 0) c143022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143022));
	wire w154022;
	repeater #(1, 1'b0, 0, 0) c154022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154022));
	wire w140023;

	wire w141023;

	wire w144023;
	repeater #(1, 1'b0, 0, 0) c144023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144023));
	wire w146023;
	repeater #(4, 1'b0, 0, 0) c146023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146023));
	wire w148023;

	wire w149023;

	wire w154023;
	repeater #(4, 1'b0, 0, 0) c154023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154023));
	wire w156023;

	wire w157023;

	wire w159023;
	repeater #(2, 1'b1, 0, 0) c159023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159023));
	wire w146024;
	repeater #(1, 1'b0, 0, 0) c146024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146024));
	wire w159024;
	repeater #(1, 1'b1, 0, 0) c159024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159024));
	wire w143025;
	repeater #(2, 1'b0, 0, 0) c143025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143025));
	wire w159025;
	repeater #(2, 1'b1, 0, 0) c159025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159025));
	wire w143026;
	repeater #(3, 1'b0, 0, 0) c143026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143026));
	wire w151026;
	repeater #(1, 1'b0, 0, 0) c151026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151026));
	wire w152026;
	repeater #(1, 1'b0, 0, 0) c152026 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152026));
	wire w151027;
	repeater #(4, 1'b0, 0, 0) c151027 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151027));
	wire w138028;

	wire w139028;

	wire w142028;
	repeater #(1, 1'b0, 0, 0) c142028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142028));
	wire w143028;

	wire w146028;

	wire w147028;

	wire w150028;
	repeater #(1, 1'b1, 0, 0) c150028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150028));
	wire w151028;

	wire w154028;

	wire w155028;

	wire w158028;
	repeater #(1, 1'b1, 0, 0) c158028 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158028));
	wire w159028;

	wire w152030;
	torch #(1'b0) c152030 (.i_clk(tick), .i_in(), .o_out(w152030));
	wire w138032;
	repeater #(1, 1'b1, 0, 0) c138032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138032));
	wire w139032;

	wire w142032;
	repeater #(1, 1'b1, 0, 0) c142032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142032));
	wire w143032;

	wire w146032;
	repeater #(1, 1'b1, 0, 0) c146032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146032));
	wire w147032;

	wire w150032;
	repeater #(1, 1'b1, 0, 0) c150032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150032));
	wire w151032;

	wire w154032;
	repeater #(1, 1'b1, 0, 0) c154032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154032));
	wire w155032;

	wire w158032;
	repeater #(1, 1'b1, 0, 0) c158032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158032));
	wire w159032;

	wire w162032;
	repeater #(1, 1'b1, 0, 0) c162032 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162032));
	wire w163032;

	wire w138036;
	repeater #(1, 1'b1, 0, 0) c138036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138036));
	wire w146036;
	repeater #(1, 1'b1, 0, 0) c146036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146036));
	wire w154036;
	repeater #(1, 1'b1, 0, 0) c154036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154036));
	wire w162036;
	repeater #(4, 1'b1, 0, 0) c162036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162036));
	wire w138037;
	repeater #(4, 1'b1, 0, 0) c138037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138037));
	wire w140037;

	wire w141037;

	wire w143037;
	repeater #(2, 1'b1, 0, 0) c143037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143037));
	wire w146037;
	repeater #(4, 1'b1, 0, 0) c146037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146037));
	wire w148037;

	wire w149037;

	wire w151037;
	repeater #(2, 1'b1, 0, 0) c151037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151037));
	wire w154037;
	repeater #(4, 1'b1, 0, 0) c154037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154037));
	wire w156037;

	wire w157037;

	wire w159037;
	repeater #(2, 1'b1, 0, 0) c159037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159037));
	wire w143038;
	repeater #(1, 1'b1, 0, 0) c143038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143038));
	wire w151038;
	repeater #(1, 1'b1, 0, 0) c151038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151038));
	wire w159038;
	repeater #(1, 1'b1, 0, 0) c159038 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159038));
	wire w143039;
	repeater #(2, 1'b1, 0, 0) c143039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143039));
	wire w151039;
	repeater #(2, 1'b1, 0, 0) c151039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151039));
	wire w159039;
	repeater #(2, 1'b1, 0, 0) c159039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159039));
	wire w162040;
	repeater #(2, 1'b1, 0, 0) c162040 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162040));
	wire w138042;

	wire w139042;

	wire w142042;
	repeater #(1, 1'b0, 0, 0) c142042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142042));
	wire w143042;

	wire w146042;

	wire w147042;

	wire w150042;
	repeater #(1, 1'b0, 0, 0) c150042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150042));
	wire w151042;

	wire w154042;

	wire w155042;

	wire w158042;
	repeater #(1, 1'b0, 0, 0) c158042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158042));
	wire w159042;

	wire w138046;
	repeater #(1, 1'b1, 0, 0) c138046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138046));
	wire w143046;
	repeater #(1, 1'b1, 0, 0) c143046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143046));
	wire w154046;
	repeater #(1, 1'b1, 0, 0) c154046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154046));
	wire w140047;

	wire w141047;

	wire w144047;
	repeater #(1, 1'b1, 0, 0) c144047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144047));
	wire w146047;
	repeater #(4, 1'b1, 0, 0) c146047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146047));
	wire w148047;

	wire w149047;

	wire w154047;
	repeater #(4, 1'b1, 0, 0) c154047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154047));
	wire w156047;

	wire w157047;

	wire w159047;
	repeater #(2, 1'b1, 0, 0) c159047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159047));
	wire w146048;
	repeater #(1, 1'b1, 0, 0) c146048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146048));
	wire w159048;
	repeater #(1, 1'b1, 0, 0) c159048 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159048));
	wire w143049;
	repeater #(2, 1'b1, 0, 0) c143049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143049));
	wire w159049;
	repeater #(2, 1'b1, 0, 0) c159049 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159049));
	wire w143050;
	repeater #(3, 1'b1, 0, 0) c143050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143050));
	wire w151050;
	repeater #(1, 1'b1, 0, 0) c151050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151050));
	wire w152050;
	repeater #(1, 1'b1, 0, 0) c152050 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152050));
	wire w151051;
	repeater #(4, 1'b1, 0, 0) c151051 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151051));
	wire w138052;

	wire w139052;

	wire w142052;
	repeater #(1, 1'b0, 0, 0) c142052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142052));
	wire w143052;

	wire w146052;

	wire w147052;

	wire w150052;
	repeater #(1, 1'b0, 0, 0) c150052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150052));
	wire w151052;

	wire w154052;

	wire w155052;

	wire w158052;
	repeater #(1, 1'b0, 0, 0) c158052 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158052));
	wire w159052;

	wire w152054;
	torch #(1'b1) c152054 (.i_clk(tick), .i_in(), .o_out(w152054));
	wire w138056;
	repeater #(1, 1'b0, 0, 0) c138056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138056));
	wire w139056;

	wire w142056;
	repeater #(1, 1'b0, 0, 0) c142056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142056));
	wire w143056;

	wire w146056;
	repeater #(1, 1'b0, 0, 0) c146056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146056));
	wire w147056;

	wire w150056;
	repeater #(1, 1'b0, 0, 0) c150056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150056));
	wire w151056;

	wire w154056;
	repeater #(1, 1'b0, 0, 0) c154056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154056));
	wire w155056;

	wire w158056;
	repeater #(1, 1'b0, 0, 0) c158056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158056));
	wire w159056;

	wire w162056;
	repeater #(1, 1'b0, 0, 0) c162056 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162056));
	wire w163056;

	wire w138060;
	repeater #(1, 1'b0, 0, 0) c138060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138060));
	wire w146060;
	repeater #(1, 1'b0, 0, 0) c146060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146060));
	wire w154060;
	repeater #(1, 1'b0, 0, 0) c154060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154060));
	wire w162060;
	repeater #(4, 1'b0, 0, 0) c162060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162060));
	wire w138061;
	repeater #(4, 1'b0, 0, 0) c138061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138061));
	wire w140061;

	wire w141061;

	wire w143061;
	repeater #(2, 1'b0, 0, 0) c143061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143061));
	wire w146061;
	repeater #(4, 1'b0, 0, 0) c146061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146061));
	wire w148061;

	wire w149061;

	wire w151061;
	repeater #(2, 1'b0, 0, 0) c151061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151061));
	wire w154061;
	repeater #(4, 1'b0, 0, 0) c154061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154061));
	wire w156061;

	wire w157061;

	wire w159061;
	repeater #(2, 1'b0, 0, 0) c159061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159061));
	wire w143062;
	repeater #(1, 1'b0, 0, 0) c143062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143062));
	wire w151062;
	repeater #(1, 1'b0, 0, 0) c151062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151062));
	wire w159062;
	repeater #(1, 1'b0, 0, 0) c159062 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159062));
	wire w143063;
	repeater #(2, 1'b0, 0, 0) c143063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143063));
	wire w151063;
	repeater #(2, 1'b0, 0, 0) c151063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151063));
	wire w159063;
	repeater #(2, 1'b0, 0, 0) c159063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159063));
	wire w162064;
	repeater #(2, 1'b0, 0, 0) c162064 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w162064));
	wire w138066;

	wire w139066;

	wire w142066;
	repeater #(1, 1'b0, 0, 0) c142066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142066));
	wire w143066;

	wire w146066;

	wire w147066;

	wire w150066;
	repeater #(1, 1'b0, 0, 0) c150066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150066));
	wire w151066;

	wire w154066;

	wire w155066;

	wire w158066;
	repeater #(1, 1'b0, 0, 0) c158066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158066));
	wire w159066;

	wire w138070;
	repeater #(1, 1'b0, 0, 0) c138070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138070));
	wire w143070;
	repeater #(1, 1'b0, 0, 0) c143070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143070));
	wire w154070;
	repeater #(1, 1'b0, 0, 0) c154070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154070));
	wire w140071;

	wire w141071;

	wire w144071;
	repeater #(1, 1'b0, 0, 0) c144071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w144071));
	wire w146071;
	repeater #(4, 1'b0, 0, 0) c146071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146071));
	wire w148071;

	wire w149071;

	wire w154071;
	repeater #(4, 1'b0, 0, 0) c154071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w154071));
	wire w156071;

	wire w157071;

	wire w159071;
	repeater #(2, 1'b0, 0, 0) c159071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159071));
	wire w146072;
	repeater #(1, 1'b0, 0, 0) c146072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146072));
	wire w159072;
	repeater #(1, 1'b0, 0, 0) c159072 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159072));
	wire w143073;
	repeater #(2, 1'b0, 0, 0) c143073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143073));
	wire w159073;
	repeater #(2, 1'b0, 0, 0) c159073 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w159073));
	wire w143074;
	repeater #(3, 1'b0, 0, 0) c143074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143074));
	wire w151074;
	repeater #(1, 1'b0, 0, 0) c151074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151074));
	wire w152074;
	repeater #(1, 1'b0, 0, 0) c152074 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w152074));
	wire w151075;
	repeater #(4, 1'b0, 0, 0) c151075 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w151075));
	wire w138076;

	wire w139076;

	wire w142076;
	repeater #(1, 1'b0, 0, 0) c142076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142076));
	wire w143076;

	wire w146076;

	wire w147076;

	wire w150076;
	repeater #(1, 1'b0, 0, 0) c150076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150076));
	wire w151076;

	wire w154076;

	wire w155076;

	wire w158076;
	repeater #(1, 1'b1, 0, 0) c158076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158076));
	wire w159076;

	wire w152078;
	torch #(1'b0) c152078 (.i_clk(tick), .i_in(), .o_out(w152078));
	wire w1370130;
	repeater #(1, 1'b0, 0, 0) c1370130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370130));
	wire w1380133;
	repeater #(1, 1'b0, 0, 0) c1380133 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380133));
	wire w1000134;
	repeater #(1, 1'b1, 0, 0) c1000134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1000134));
	wire w1170134;
	repeater #(2, 1'b1, 0, 0) c1170134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1170134));
	wire w1180134;
	repeater #(1, 1'b1, 0, 0) c1180134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1180134));
	wire w1190134;

	wire w1340134;

	wire w1370134;
	repeater #(1, 1'b1, 0, 0) c1370134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1370134));
	wire w1470134;
	repeater #(1, 1'b1, 0, 0) c1470134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470134));
	wire w1520134;
	repeater #(1, 1'b1, 0, 0) c1520134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1520134));
	wire w1360135;
	repeater #(1, 1'b0, 0, 0) c1360135 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1360135));
	wire w1490135;

	wire w1500135;

	wire w1500137;
	repeater #(1, 1'b0, 0, 0) c1500137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500137));
	wire w1640137;
	repeater #(1, 1'b1, 0, 0) c1640137 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640137));
	wire w1350138;
	repeater #(1, 1'b0, 0, 0) c1350138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350138));
	wire w1640138;

	wire w1660139;
	repeater #(1, 1'b0, 0, 0) c1660139 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1660139));
	wire w1390145;
	repeater #(1, 1'b0, 0, 0) c1390145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390145));
	wire w1420145;
	repeater #(1, 1'b0, 0, 0) c1420145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420145));
	wire w1470145;
	repeater #(1, 1'b0, 0, 0) c1470145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470145));
	wire w1500145;
	repeater #(1, 1'b0, 0, 0) c1500145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500145));
	wire w1550145;
	repeater #(1, 1'b0, 0, 0) c1550145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550145));
	wire w1580145;
	repeater #(1, 1'b0, 0, 0) c1580145 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580145));
	wire w1380154;
	repeater #(3, 1'b0, 0, 0) c1380154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380154));
	wire w1470155;
	repeater #(1, 1'b0, 0, 0) c1470155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470155));
	wire w1500155;
	repeater #(1, 1'b0, 0, 0) c1500155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500155));
	wire w1550155;
	repeater #(1, 1'b0, 0, 0) c1550155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550155));
	wire w1580155;
	repeater #(1, 1'b0, 0, 0) c1580155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580155));
	wire w1660155;
	repeater #(1, 1'b0, 0, 0) c1660155 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1660155));
	wire w1640159;
	repeater #(1, 1'b1, 0, 0) c1640159 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640159));
	wire w1640161;
	repeater #(1, 1'b1, 0, 0) c1640161 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1640161));
	wire w1640162;

	wire w1660163;
	repeater #(1, 1'b0, 0, 0) c1660163 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1660163));
	wire w1390169;
	repeater #(1, 1'b1, 0, 0) c1390169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1390169));
	wire w1420169;
	repeater #(1, 1'b1, 0, 0) c1420169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420169));
	wire w1470169;
	repeater #(1, 1'b1, 0, 0) c1470169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1470169));
	wire w1500169;
	repeater #(1, 1'b1, 0, 0) c1500169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1500169));
	wire w1550169;
	repeater #(1, 1'b1, 0, 0) c1550169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1550169));
	wire w1580169;
	repeater #(1, 1'b1, 0, 0) c1580169 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1580169));
	wire w1380178;
	repeater #(3, 1'b1, 0, 0) c1380178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380178));
	wire w14710;
	repeater #(1, 1'b1, 0, 0) c14710 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w14710));
	wire w15010;
	repeater #(1, 1'b1, 0, 0) c15010 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15010));
	wire w15510;
	repeater #(1, 1'b1, 0, 0) c15510 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15510));
	wire w15810;
	repeater #(1, 1'b1, 0, 0) c15810 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w15810));
	wire w16610;
	repeater #(1, 1'b0, 0, 0) c16610 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16610));
	wire w16414;
	repeater #(1, 1'b1, 0, 0) c16414 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16414));
	wire w16416;
	repeater #(1, 1'b1, 0, 0) c16416 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16416));
	wire w16417;

	wire w16618;
	repeater #(1, 1'b0, 0, 0) c16618 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w16618));
	wire w139114;
	repeater #(1, 1'b0, 0, 0) c139114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139114));
	wire w142114;
	repeater #(1, 1'b0, 0, 0) c142114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142114));
	wire w147114;
	repeater #(1, 1'b0, 0, 0) c147114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147114));
	wire w150114;
	repeater #(1, 1'b0, 0, 0) c150114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150114));
	wire w155114;
	repeater #(1, 1'b1, 0, 0) c155114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155114));
	wire w158114;
	repeater #(1, 1'b0, 0, 0) c158114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158114));
	wire w138123;
	repeater #(3, 1'b0, 0, 0) c138123 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138123));
	wire w147124;
	repeater #(1, 1'b0, 0, 0) c147124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147124));
	wire w150124;
	repeater #(1, 1'b0, 0, 0) c150124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150124));
	wire w155124;
	repeater #(1, 1'b1, 0, 0) c155124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155124));
	wire w158124;
	repeater #(1, 1'b0, 0, 0) c158124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158124));
	wire w166124;
	repeater #(1, 1'b0, 0, 0) c166124 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166124));
	wire w164128;
	repeater #(1, 1'b1, 0, 0) c164128 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164128));
	wire w164130;
	repeater #(1, 1'b1, 0, 0) c164130 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164130));
	wire w164131;

	wire w166132;
	repeater #(1, 1'b0, 0, 0) c166132 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166132));
	wire w139138;
	repeater #(1, 1'b1, 0, 0) c139138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139138));
	wire w142138;
	repeater #(1, 1'b1, 0, 0) c142138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142138));
	wire w147138;
	repeater #(1, 1'b1, 0, 0) c147138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147138));
	wire w150138;
	repeater #(1, 1'b1, 0, 0) c150138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150138));
	wire w155138;
	repeater #(1, 1'b1, 0, 0) c155138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155138));
	wire w158138;
	repeater #(1, 1'b1, 0, 0) c158138 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158138));
	wire w138147;
	repeater #(3, 1'b1, 0, 0) c138147 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138147));
	wire w147148;
	repeater #(1, 1'b1, 0, 0) c147148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147148));
	wire w150148;
	repeater #(1, 1'b1, 0, 0) c150148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150148));
	wire w155148;
	repeater #(1, 1'b1, 0, 0) c155148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155148));
	wire w158148;
	repeater #(1, 1'b1, 0, 0) c158148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158148));
	wire w166148;
	repeater #(1, 1'b0, 0, 0) c166148 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166148));
	wire w164152;
	repeater #(1, 1'b1, 0, 0) c164152 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164152));
	wire w164154;
	repeater #(1, 1'b1, 0, 0) c164154 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164154));
	wire w164155;

	wire w166156;
	repeater #(1, 1'b0, 0, 0) c166156 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166156));
	wire w139162;
	repeater #(1, 1'b0, 0, 0) c139162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w139162));
	wire w142162;
	repeater #(1, 1'b0, 0, 0) c142162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142162));
	wire w147162;
	repeater #(1, 1'b0, 0, 0) c147162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147162));
	wire w150162;
	repeater #(1, 1'b0, 0, 0) c150162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150162));
	wire w155162;
	repeater #(1, 1'b0, 0, 0) c155162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155162));
	wire w158162;
	repeater #(1, 1'b0, 0, 0) c158162 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158162));
	wire w138171;
	repeater #(3, 1'b0, 0, 0) c138171 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138171));
	wire w147172;
	repeater #(1, 1'b0, 0, 0) c147172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w147172));
	wire w150172;
	repeater #(1, 1'b0, 0, 0) c150172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w150172));
	wire w155172;
	repeater #(1, 1'b0, 0, 0) c155172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w155172));
	wire w158172;
	repeater #(1, 1'b0, 0, 0) c158172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w158172));
	wire w166172;
	repeater #(1, 1'b0, 0, 0) c166172 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w166172));
	wire w164174;
	torch #(1'b0) c164174 (.i_clk(tick), .i_in(), .o_out(w164174));
	wire w164176;
	repeater #(1, 1'b0, 0, 0) c164176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164176));
	wire w168177;
	repeater #(1, 1'b0, 0, 0) c168177 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w168177));
	wire w164178;
	repeater #(1, 1'b0, 0, 0) c164178 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w164178));
	wire w164179;

	wire w169179;

	wire w172179;
	assign outputs[125] = ();
	wire w169180;

	wire w167181;
	repeater #(1, 1'b0, 0, 0) c167181 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w167181));
	wire w122012;
	repeater #(1, 1'b0, 0, 0) c122012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122012));
	wire w127012;
	repeater #(1, 1'b0, 0, 0) c127012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127012));
	wire w130012;
	repeater #(1, 1'b1, 0, 0) c130012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130012));
	wire w135012;
	repeater #(1, 1'b0, 0, 0) c135012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135012));
	wire w138012;
	repeater #(1, 1'b0, 0, 0) c138012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138012));
	wire w143012;
	repeater #(1, 1'b0, 0, 0) c143012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143012));
	wire w146012;
	repeater #(1, 1'b0, 0, 0) c146012 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146012));
	wire w122013;

	wire w123013;

	wire w126013;
	repeater #(1, 1'b0, 0, 0) c126013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126013));
	wire w127013;

	wire w130013;

	wire w131013;

	wire w134013;
	repeater #(1, 1'b1, 0, 0) c134013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134013));
	wire w135013;

	wire w138013;

	wire w139013;

	wire w142013;
	repeater #(1, 1'b1, 0, 0) c142013 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142013));
	wire w143013;

	wire w146013;

	wire w124017;
	repeater #(1, 1'b0, 0, 0) c124017 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124017));
	wire w123018;
	repeater #(1, 1'b0, 0, 0) c123018 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123018));
	wire w122022;
	repeater #(1, 1'b0, 0, 0) c122022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122022));
	wire w127022;
	repeater #(1, 1'b1, 0, 0) c127022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127022));
	wire w130022;
	repeater #(1, 1'b1, 0, 0) c130022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130022));
	wire w135022;
	repeater #(1, 1'b0, 0, 0) c135022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135022));
	wire w138022;
	repeater #(1, 1'b0, 0, 0) c138022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138022));
	wire w143022;
	repeater #(1, 1'b0, 0, 0) c143022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143022));
	wire w122023;

	wire w123023;

	wire w126023;
	repeater #(1, 1'b0, 0, 0) c126023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126023));
	wire w127023;

	wire w130023;

	wire w131023;

	wire w134023;
	repeater #(1, 1'b1, 0, 0) c134023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134023));
	wire w135023;

	wire w138023;

	wire w139023;

	wire w142023;
	repeater #(1, 1'b1, 0, 0) c142023 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142023));
	wire w143023;

	wire w122036;
	repeater #(1, 1'b0, 0, 0) c122036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122036));
	wire w127036;
	repeater #(1, 1'b0, 0, 0) c127036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127036));
	wire w130036;
	repeater #(1, 1'b0, 0, 0) c130036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130036));
	wire w135036;
	repeater #(1, 1'b1, 0, 0) c135036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135036));
	wire w138036;
	repeater #(1, 1'b0, 0, 0) c138036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138036));
	wire w143036;
	repeater #(1, 1'b0, 0, 0) c143036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143036));
	wire w146036;
	repeater #(1, 1'b0, 0, 0) c146036 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146036));
	wire w122037;

	wire w123037;

	wire w126037;
	repeater #(1, 1'b1, 0, 0) c126037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126037));
	wire w127037;

	wire w130037;

	wire w131037;

	wire w134037;
	repeater #(1, 1'b0, 0, 0) c134037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134037));
	wire w135037;

	wire w138037;

	wire w139037;

	wire w142037;
	repeater #(1, 1'b1, 0, 0) c142037 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142037));
	wire w143037;

	wire w146037;

	wire w124041;
	repeater #(1, 1'b1, 0, 0) c124041 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124041));
	wire w123042;
	repeater #(1, 1'b1, 0, 0) c123042 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123042));
	wire w122046;
	repeater #(1, 1'b0, 0, 0) c122046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122046));
	wire w127046;
	repeater #(1, 1'b1, 0, 0) c127046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127046));
	wire w130046;
	repeater #(1, 1'b1, 0, 0) c130046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130046));
	wire w135046;
	repeater #(1, 1'b0, 0, 0) c135046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135046));
	wire w138046;
	repeater #(1, 1'b0, 0, 0) c138046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138046));
	wire w143046;
	repeater #(1, 1'b0, 0, 0) c143046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143046));
	wire w122047;

	wire w123047;

	wire w126047;
	repeater #(1, 1'b0, 0, 0) c126047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126047));
	wire w127047;

	wire w130047;

	wire w131047;

	wire w134047;
	repeater #(1, 1'b1, 0, 0) c134047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134047));
	wire w135047;

	wire w138047;

	wire w139047;

	wire w142047;
	repeater #(1, 1'b1, 0, 0) c142047 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142047));
	wire w143047;

	wire w122060;
	repeater #(1, 1'b0, 0, 0) c122060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122060));
	wire w127060;
	repeater #(1, 1'b0, 0, 0) c127060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127060));
	wire w130060;
	repeater #(1, 1'b0, 0, 0) c130060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130060));
	wire w135060;
	repeater #(1, 1'b1, 0, 0) c135060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135060));
	wire w138060;
	repeater #(1, 1'b0, 0, 0) c138060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138060));
	wire w143060;
	repeater #(1, 1'b0, 0, 0) c143060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143060));
	wire w146060;
	repeater #(1, 1'b0, 0, 0) c146060 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146060));
	wire w122061;

	wire w123061;

	wire w126061;
	repeater #(1, 1'b0, 0, 0) c126061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126061));
	wire w127061;

	wire w130061;

	wire w131061;

	wire w134061;
	repeater #(1, 1'b0, 0, 0) c134061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134061));
	wire w135061;

	wire w138061;

	wire w139061;

	wire w142061;
	repeater #(1, 1'b1, 0, 0) c142061 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142061));
	wire w143061;

	wire w146061;

	wire w124065;
	repeater #(1, 1'b0, 0, 0) c124065 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124065));
	wire w123066;
	repeater #(1, 1'b0, 0, 0) c123066 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123066));
	wire w122070;
	repeater #(1, 1'b0, 0, 0) c122070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122070));
	wire w127070;
	repeater #(1, 1'b1, 0, 0) c127070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127070));
	wire w130070;
	repeater #(1, 1'b1, 0, 0) c130070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130070));
	wire w135070;
	repeater #(1, 1'b0, 0, 0) c135070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135070));
	wire w138070;
	repeater #(1, 1'b0, 0, 0) c138070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138070));
	wire w143070;
	repeater #(1, 1'b0, 0, 0) c143070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143070));
	wire w122071;

	wire w123071;

	wire w126071;
	repeater #(1, 1'b0, 0, 0) c126071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126071));
	wire w127071;

	wire w130071;

	wire w131071;

	wire w134071;
	repeater #(1, 1'b1, 0, 0) c134071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134071));
	wire w135071;

	wire w138071;

	wire w139071;

	wire w142071;
	repeater #(1, 1'b1, 0, 0) c142071 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142071));
	wire w143071;

	wire w122084;
	repeater #(1, 1'b0, 0, 0) c122084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122084));
	wire w127084;
	repeater #(1, 1'b0, 0, 0) c127084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127084));
	wire w130084;
	repeater #(1, 1'b0, 0, 0) c130084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130084));
	wire w135084;
	repeater #(1, 1'b0, 0, 0) c135084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135084));
	wire w138084;
	repeater #(1, 1'b0, 0, 0) c138084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138084));
	wire w143084;
	repeater #(1, 1'b0, 0, 0) c143084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143084));
	wire w146084;
	repeater #(1, 1'b1, 0, 0) c146084 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w146084));
	wire w122085;

	wire w123085;

	wire w126085;
	repeater #(1, 1'b0, 0, 0) c126085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126085));
	wire w127085;

	wire w130085;

	wire w131085;

	wire w134085;
	repeater #(1, 1'b0, 0, 0) c134085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134085));
	wire w135085;

	wire w138085;

	wire w139085;

	wire w142085;
	repeater #(1, 1'b0, 0, 0) c142085 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142085));
	wire w143085;

	wire w146085;

	wire w124089;
	repeater #(1, 1'b1, 0, 0) c124089 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w124089));
	wire w123090;
	repeater #(1, 1'b1, 0, 0) c123090 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w123090));
	wire w122094;
	repeater #(1, 1'b0, 0, 0) c122094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w122094));
	wire w127094;
	repeater #(1, 1'b0, 0, 0) c127094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w127094));
	wire w130094;
	repeater #(1, 1'b0, 0, 0) c130094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w130094));
	wire w135094;
	repeater #(1, 1'b1, 0, 0) c135094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w135094));
	wire w138094;
	repeater #(1, 1'b0, 0, 0) c138094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w138094));
	wire w143094;
	repeater #(1, 1'b1, 0, 0) c143094 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w143094));
	wire w122095;

	wire w123095;

	wire w126095;
	repeater #(1, 1'b0, 0, 0) c126095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w126095));
	wire w127095;

	wire w130095;

	wire w131095;

	wire w134095;
	repeater #(1, 1'b0, 0, 0) c134095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w134095));
	wire w135095;

	wire w138095;

	wire w139095;

	wire w142095;
	repeater #(1, 1'b0, 0, 0) c142095 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w142095));
	wire w143095;

	wire w1220108;
	repeater #(1, 1'b0, 0, 0) c1220108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1220108));
	wire w1270108;
	repeater #(1, 1'b0, 0, 0) c1270108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1270108));
	wire w1300108;
	repeater #(1, 1'b0, 0, 0) c1300108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1300108));
	wire w1350108;
	repeater #(1, 1'b0, 0, 0) c1350108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350108));
	wire w1380108;
	repeater #(1, 1'b0, 0, 0) c1380108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380108));
	wire w1430108;
	repeater #(1, 1'b1, 0, 0) c1430108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1430108));
	wire w1460108;
	repeater #(1, 1'b0, 0, 0) c1460108 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1460108));
	wire w1220109;

	wire w1230109;

	wire w1260109;
	repeater #(1, 1'b0, 0, 0) c1260109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1260109));
	wire w1270109;

	wire w1300109;

	wire w1310109;

	wire w1340109;
	repeater #(1, 1'b0, 0, 0) c1340109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340109));
	wire w1350109;

	wire w1380109;

	wire w1390109;

	wire w1420109;
	repeater #(1, 1'b0, 0, 0) c1420109 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420109));
	wire w1430109;

	wire w1460109;

	wire w1240113;
	repeater #(1, 1'b0, 0, 0) c1240113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1240113));
	wire w1230114;
	repeater #(1, 1'b0, 0, 0) c1230114 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1230114));
	wire w1220118;
	repeater #(1, 1'b0, 0, 0) c1220118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1220118));
	wire w1270118;
	repeater #(1, 1'b0, 0, 0) c1270118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1270118));
	wire w1300118;
	repeater #(1, 1'b0, 0, 0) c1300118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1300118));
	wire w1350118;
	repeater #(1, 1'b1, 0, 0) c1350118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1350118));
	wire w1380118;
	repeater #(1, 1'b1, 0, 0) c1380118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1380118));
	wire w1430118;
	repeater #(1, 1'b0, 0, 0) c1430118 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1430118));
	wire w1220119;

	wire w1230119;

	wire w1260119;
	repeater #(1, 1'b0, 0, 0) c1260119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1260119));
	wire w1270119;

	wire w1300119;

	wire w1310119;

	wire w1340119;
	repeater #(1, 1'b0, 0, 0) c1340119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1340119));
	wire w1350119;

	wire w1380119;

	wire w1390119;

	wire w1420119;
	repeater #(1, 1'b1, 0, 0) c1420119 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1420119));
	wire w1430119;

	wire w106162;

	wire w110162;

	wire w114162;

	wire w118162;

	wire w122162;

	wire w126162;

	wire w130162;

	wire w105164;
	repeater #(1, 1'b1, 0, 0) c105164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105164));
	wire w113164;
	repeater #(1, 1'b1, 0, 0) c113164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113164));
	wire w121164;
	repeater #(2, 1'b1, 0, 0) c121164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121164));
	wire w129164;
	repeater #(2, 1'b1, 0, 0) c129164 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w129164));
	wire w120165;
	repeater #(1, 1'b1, 0, 0) c120165 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120165));
	wire w106186;

	wire w110186;

	wire w114186;

	wire w118186;

	wire w122186;

	wire w126186;

	wire w130186;

	wire w105188;
	repeater #(1, 1'b1, 0, 0) c105188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105188));
	wire w113188;
	repeater #(1, 1'b1, 0, 0) c113188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113188));
	wire w121188;
	repeater #(2, 1'b1, 0, 0) c121188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w121188));
	wire w129188;
	repeater #(2, 1'b1, 0, 0) c129188 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w129188));
	wire w120189;
	repeater #(1, 1'b1, 0, 0) c120189 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w120189));
	wire w1061110;

	wire w1101110;

	wire w1141110;

	wire w1181110;

	wire w1221110;

	wire w1261110;

	wire w1301110;

	wire w1051112;
	repeater #(1, 1'b1, 0, 0) c1051112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1051112));
	wire w1131112;
	repeater #(1, 1'b1, 0, 0) c1131112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1131112));
	wire w1211112;
	repeater #(2, 1'b1, 0, 0) c1211112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1211112));
	wire w1291112;
	repeater #(2, 1'b1, 0, 0) c1291112 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1291112));
	wire w1201113;
	repeater #(1, 1'b1, 0, 0) c1201113 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1201113));
	wire w1061134;

	wire w1101134;

	wire w1141134;

	wire w1181134;

	wire w1221134;

	wire w1261134;

	wire w1301134;

	wire w8900;
	repeater #(1, 1'b1, 0, 0) c8900 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w8900));
	wire w9700;
	repeater #(1, 1'b1, 0, 0) c9700 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w9700));
	wire w10500;
	repeater #(2, 1'b1, 0, 0) c10500 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10500));
	wire w11300;
	repeater #(2, 1'b1, 0, 0) c11300 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w11300));
	wire w10401;
	repeater #(1, 1'b1, 0, 0) c10401 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w10401));
	wire w90022;

	wire w94022;

	wire w98022;

	wire w102022;

	wire w106022;

	wire w110022;

	wire w114022;

	wire w89024;
	repeater #(1, 1'b1, 0, 0) c89024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w89024));
	wire w97024;
	repeater #(1, 1'b1, 0, 0) c97024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w97024));
	wire w105024;
	repeater #(2, 1'b1, 0, 0) c105024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w105024));
	wire w113024;
	repeater #(2, 1'b1, 0, 0) c113024 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w113024));
	wire w104025;
	repeater #(1, 1'b1, 0, 0) c104025 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w104025));
	wire w901110;
	repeater #(1, 1'b0, 0, 0) c901110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901110));
	wire w941110;
	repeater #(1, 1'b0, 0, 0) c941110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941110));
	wire w981110;
	repeater #(1, 1'b0, 0, 0) c981110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981110));
	wire w1021110;
	repeater #(1, 1'b0, 0, 0) c1021110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1021110));
	wire w1061110;
	repeater #(1, 1'b0, 0, 0) c1061110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061110));
	wire w1101110;
	repeater #(1, 1'b0, 0, 0) c1101110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101110));
	wire w1141110;
	repeater #(1, 1'b0, 0, 0) c1141110 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1141110));
	wire w901127;
	repeater #(1, 1'b0, 0, 0) c901127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901127));
	wire w941127;
	repeater #(1, 1'b0, 0, 0) c941127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941127));
	wire w981127;
	repeater #(1, 1'b0, 0, 0) c981127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981127));
	wire w1021127;
	repeater #(1, 1'b0, 0, 0) c1021127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1021127));
	wire w1061127;
	repeater #(1, 1'b0, 0, 0) c1061127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061127));
	wire w1101127;
	repeater #(1, 1'b0, 0, 0) c1101127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101127));
	wire w1141127;
	repeater #(1, 1'b0, 0, 0) c1141127 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1141127));
	wire w901134;
	repeater #(1, 1'b0, 0, 0) c901134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w901134));
	wire w941134;
	repeater #(1, 1'b0, 0, 0) c941134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w941134));
	wire w981134;
	repeater #(1, 1'b0, 0, 0) c981134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w981134));
	wire w1021134;
	repeater #(1, 1'b0, 0, 0) c1021134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1021134));
	wire w1061134;
	repeater #(1, 1'b0, 0, 0) c1061134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1061134));
	wire w1101134;
	repeater #(1, 1'b0, 0, 0) c1101134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1101134));
	wire w1141134;
	repeater #(1, 1'b0, 0, 0) c1141134 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w1141134));
	wire w74015;
	repeater #(1, 1'b0, 0, 0) c74015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74015));
	wire w78015;
	repeater #(1, 1'b0, 0, 0) c78015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78015));
	wire w82015;
	repeater #(1, 1'b0, 0, 0) c82015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82015));
	wire w86015;
	repeater #(1, 1'b0, 0, 0) c86015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86015));
	wire w90015;
	repeater #(1, 1'b0, 0, 0) c90015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90015));
	wire w94015;
	repeater #(1, 1'b0, 0, 0) c94015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94015));
	wire w98015;
	repeater #(1, 1'b0, 0, 0) c98015 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98015));
	wire w74022;
	repeater #(1, 1'b0, 0, 0) c74022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74022));
	wire w78022;
	repeater #(1, 1'b0, 0, 0) c78022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78022));
	wire w82022;
	repeater #(1, 1'b0, 0, 0) c82022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82022));
	wire w86022;
	repeater #(1, 1'b0, 0, 0) c86022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86022));
	wire w90022;
	repeater #(1, 1'b0, 0, 0) c90022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90022));
	wire w94022;
	repeater #(1, 1'b0, 0, 0) c94022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94022));
	wire w98022;
	repeater #(1, 1'b0, 0, 0) c98022 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98022));
	wire w74039;
	repeater #(1, 1'b0, 0, 0) c74039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74039));
	wire w78039;
	repeater #(1, 1'b0, 0, 0) c78039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78039));
	wire w82039;
	repeater #(1, 1'b0, 0, 0) c82039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82039));
	wire w86039;
	repeater #(1, 1'b0, 0, 0) c86039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86039));
	wire w90039;
	repeater #(1, 1'b0, 0, 0) c90039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90039));
	wire w94039;
	repeater #(1, 1'b0, 0, 0) c94039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94039));
	wire w98039;
	repeater #(1, 1'b0, 0, 0) c98039 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98039));
	wire w74046;
	repeater #(1, 1'b0, 0, 0) c74046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74046));
	wire w78046;
	repeater #(1, 1'b0, 0, 0) c78046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78046));
	wire w82046;
	repeater #(1, 1'b0, 0, 0) c82046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82046));
	wire w86046;
	repeater #(1, 1'b0, 0, 0) c86046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86046));
	wire w90046;
	repeater #(1, 1'b0, 0, 0) c90046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90046));
	wire w94046;
	repeater #(1, 1'b0, 0, 0) c94046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94046));
	wire w98046;
	repeater #(1, 1'b0, 0, 0) c98046 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98046));
	wire w74063;
	repeater #(1, 1'b0, 0, 0) c74063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74063));
	wire w78063;
	repeater #(1, 1'b0, 0, 0) c78063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78063));
	wire w82063;
	repeater #(1, 1'b0, 0, 0) c82063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82063));
	wire w86063;
	repeater #(1, 1'b0, 0, 0) c86063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86063));
	wire w90063;
	repeater #(1, 1'b0, 0, 0) c90063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90063));
	wire w94063;
	repeater #(1, 1'b0, 0, 0) c94063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94063));
	wire w98063;
	repeater #(1, 1'b0, 0, 0) c98063 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98063));
	wire w74070;
	repeater #(1, 1'b0, 0, 0) c74070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w74070));
	wire w78070;
	repeater #(1, 1'b0, 0, 0) c78070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w78070));
	wire w82070;
	repeater #(1, 1'b0, 0, 0) c82070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w82070));
	wire w86070;
	repeater #(1, 1'b0, 0, 0) c86070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w86070));
	wire w90070;
	repeater #(1, 1'b0, 0, 0) c90070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w90070));
	wire w94070;
	repeater #(1, 1'b0, 0, 0) c94070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w94070));
	wire w98070;
	repeater #(1, 1'b0, 0, 0) c98070 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w98070));
	wire w74076;

	wire w75076;
	repeater #(1, 1'b1, 0, 0) c75076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w75076));
	wire w78076;

	wire w79076;
	repeater #(1, 1'b1, 0, 0) c79076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w79076));
	wire w82076;

	wire w83076;
	repeater #(1, 1'b1, 0, 0) c83076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w83076));
	wire w86076;

	wire w87076;
	repeater #(1, 1'b1, 0, 0) c87076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w87076));
	wire w90076;

	wire w91076;
	repeater #(1, 1'b1, 0, 0) c91076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w91076));
	wire w94076;

	wire w95076;
	repeater #(1, 1'b1, 0, 0) c95076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w95076));
	wire w98076;

	wire w99076;
	repeater #(1, 1'b1, 0, 0) c99076 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w99076));
	wire w101076;
	assign w101076 = inputs[21];
	wire w85176;
	repeater #(1, 1'b1, 0, 0) c85176 (.i_clk(tick), .i_in(), .i_lock(), .o_out(w85176));
endmodule