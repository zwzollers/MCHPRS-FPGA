module redstone (tick, inputs, outputs);
	input tick;
	input [num_inputs-1:0] inputs;
	output [num_outputs:0] outputs;

parameter num_outputs = 1, num_inputs = 1;

	wire w112;
	assign w112 = inputs[0];
	wire w121;
	torch #(1'b0) c121 (.i_clk(tick), .i_in(w112), .o_out(w121));
	wire w132;
	torch #(1'b1) c132 (.i_clk(tick), .i_in(w121|w142), .o_out(w132));
	wire w142;
	repeater #(1, 1'b0, 0, 0) c142 (.i_clk(tick), .i_in(w132), .i_lock(), .o_out(w142));
	wire w154;
	torch #(1'b0) c154 (.i_clk(tick), .i_in(w132), .o_out(w154));
	wire w192;
	repeater #(1, 1'b1, 0, 0) c192 (.i_clk(tick), .i_in(w154), .i_lock(), .o_out(w192));
	wire w199;
	repeater #(1, 1'b1, 0, 0) c199 (.i_clk(tick), .i_in(w154), .i_lock(), .o_out(w199));
	wire w204;
	repeater #(1, 1'b1, 1, 0) c204 (.i_clk(tick), .i_in(w192), .i_lock(), .o_out(w204));
	wire w205;
	repeater #(1, 1'b1, 0, 1) c205 (.i_clk(tick), .i_in(w206), .i_lock(w204), .o_out(w205));
	wire w206;
	repeater #(1, 1'b0, 0, 1) c206 (.i_clk(tick), .i_in(w205), .i_lock(w207), .o_out(w206));
	wire w207;
	repeater #(1, 1'b1, 1, 0) c207 (.i_clk(tick), .i_in(w199), .i_lock(), .o_out(w207));
	wire w294;
	repeater #(1, 1'b1, 0, 0) c294 (.i_clk(tick), .i_in(w205), .i_lock(), .o_out(w294));
	wire w297;
	repeater #(1, 1'b1, 0, 0) c297 (.i_clk(tick), .i_in(w205), .i_lock(), .o_out(w297));
	wire w424;
	repeater #(1, 1'b1, 1, 0) c424 (.i_clk(tick), .i_in(w192|w294), .i_lock(), .o_out(w424));
	wire w425;
	repeater #(1, 1'b1, 0, 1) c425 (.i_clk(tick), .i_in(w426), .i_lock(w424), .o_out(w425));
	wire w426;
	repeater #(1, 1'b0, 0, 1) c426 (.i_clk(tick), .i_in(w425), .i_lock(w427), .o_out(w426));
	wire w427;
	repeater #(1, 1'b1, 1, 0) c427 (.i_clk(tick), .i_in(w199|w297), .i_lock(), .o_out(w427));
	wire w514;
	repeater #(1, 1'b1, 0, 0) c514 (.i_clk(tick), .i_in(w425), .i_lock(), .o_out(w514));
	wire w517;
	repeater #(1, 1'b1, 0, 0) c517 (.i_clk(tick), .i_in(w425), .i_lock(), .o_out(w517));
	wire w644;
	repeater #(1, 1'b1, 1, 0) c644 (.i_clk(tick), .i_in(w192|w294|w514), .i_lock(), .o_out(w644));
	wire w645;
	repeater #(1, 1'b1, 0, 1) c645 (.i_clk(tick), .i_in(w646), .i_lock(w644), .o_out(w645));
	wire w646;
	repeater #(1, 1'b0, 0, 1) c646 (.i_clk(tick), .i_in(w645), .i_lock(w647), .o_out(w646));
	wire w647;
	repeater #(1, 1'b1, 1, 0) c647 (.i_clk(tick), .i_in(w199|w297|w517), .i_lock(), .o_out(w647));
	wire w734;
	repeater #(1, 1'b1, 0, 0) c734 (.i_clk(tick), .i_in(w645), .i_lock(), .o_out(w734));
	wire w737;
	repeater #(1, 1'b1, 0, 0) c737 (.i_clk(tick), .i_in(w645), .i_lock(), .o_out(w737));
	wire w864;
	repeater #(1, 1'b1, 1, 0) c864 (.i_clk(tick), .i_in(w192|w294|w514|w734), .i_lock(), .o_out(w864));
	wire w865;
	repeater #(1, 1'b1, 0, 1) c865 (.i_clk(tick), .i_in(w866), .i_lock(w864), .o_out(w865));
	wire w866;
	repeater #(1, 1'b0, 0, 1) c866 (.i_clk(tick), .i_in(w865), .i_lock(w867), .o_out(w866));
	wire w867;
	repeater #(1, 1'b1, 1, 0) c867 (.i_clk(tick), .i_in(w199|w297|w517|w737), .i_lock(), .o_out(w867));
	wire w954;
	repeater #(1, 1'b1, 0, 0) c954 (.i_clk(tick), .i_in(w865), .i_lock(), .o_out(w954));
	wire w957;
	repeater #(1, 1'b1, 0, 0) c957 (.i_clk(tick), .i_in(w865), .i_lock(), .o_out(w957));
	wire w1084;
	repeater #(1, 1'b1, 1, 0) c1084 (.i_clk(tick), .i_in(w192|w294|w514|w734|w954), .i_lock(), .o_out(w1084));
	wire w1085;
	repeater #(1, 1'b1, 0, 1) c1085 (.i_clk(tick), .i_in(w1086), .i_lock(w1084), .o_out(w1085));
	wire w1086;
	repeater #(1, 1'b0, 0, 1) c1086 (.i_clk(tick), .i_in(w1085), .i_lock(w1087), .o_out(w1086));
	wire w1087;
	repeater #(1, 1'b1, 1, 0) c1087 (.i_clk(tick), .i_in(w199|w297|w517|w737|w957), .i_lock(), .o_out(w1087));
	wire w1174;
	repeater #(1, 1'b1, 0, 0) c1174 (.i_clk(tick), .i_in(w1085), .i_lock(), .o_out(w1174));
	wire w1177;
	repeater #(1, 1'b1, 0, 0) c1177 (.i_clk(tick), .i_in(w1085), .i_lock(), .o_out(w1177));
	wire w1304;
	repeater #(1, 1'b1, 1, 0) c1304 (.i_clk(tick), .i_in(w192|w294|w514|w734|w954|w1174), .i_lock(), .o_out(w1304));
	wire w1305;
	repeater #(1, 1'b1, 0, 1) c1305 (.i_clk(tick), .i_in(w1306), .i_lock(w1304), .o_out(w1305));
	wire w1306;
	repeater #(1, 1'b0, 0, 1) c1306 (.i_clk(tick), .i_in(w1305), .i_lock(w1307), .o_out(w1306));
	wire w1307;
	repeater #(1, 1'b1, 1, 0) c1307 (.i_clk(tick), .i_in(w199|w297|w517|w737|w957|w1177), .i_lock(), .o_out(w1307));
	wire w1394;
	repeater #(1, 1'b1, 0, 0) c1394 (.i_clk(tick), .i_in(w1305), .i_lock(), .o_out(w1394));
	wire w1397;
	repeater #(1, 1'b1, 0, 0) c1397 (.i_clk(tick), .i_in(w1305), .i_lock(), .o_out(w1397));
	wire w1524;
	repeater #(1, 1'b1, 1, 0) c1524 (.i_clk(tick), .i_in(w192|w294|w514|w734|w954|w1174|w1394), .i_lock(), .o_out(w1524));
	wire w1525;
	repeater #(1, 1'b1, 0, 1) c1525 (.i_clk(tick), .i_in(w1526), .i_lock(w1524), .o_out(w1525));
	wire w1526;
	repeater #(1, 1'b0, 0, 1) c1526 (.i_clk(tick), .i_in(w1525), .i_lock(w1527), .o_out(w1526));
	wire w1527;
	repeater #(1, 1'b1, 1, 0) c1527 (.i_clk(tick), .i_in(w199|w297|w517|w737|w957|w1177|w1397), .i_lock(), .o_out(w1527));
	wire w1614;
	repeater #(1, 1'b1, 0, 0) c1614 (.i_clk(tick), .i_in(w1525), .i_lock(), .o_out(w1614));
	wire w1617;
	repeater #(1, 1'b1, 0, 0) c1617 (.i_clk(tick), .i_in(w1525), .i_lock(), .o_out(w1617));
	wire w1685;
	torch #(1'b1) c1685 (.i_clk(tick), .i_in(w1745), .o_out(w1685));
	wire w1686;
	repeater #(2, 1'b0, 0, 0) c1686 (.i_clk(tick), .i_in(w1685), .i_lock(), .o_out(w1686));
	wire w1696;
	repeater #(1, 1'b1, 0, 0) c1696 (.i_clk(tick), .i_in(w1745), .i_lock(), .o_out(w1696));
	wire w1744;
	repeater #(1, 1'b1, 1, 0) c1744 (.i_clk(tick), .i_in(w192|w294|w514|w734|w954|w1174|w1394|w1614), .i_lock(), .o_out(w1744));
	wire w1745;
	repeater #(1, 1'b1, 0, 1) c1745 (.i_clk(tick), .i_in(w1746), .i_lock(w1744), .o_out(w1745));
	wire w1746;
	repeater #(1, 1'b0, 0, 1) c1746 (.i_clk(tick), .i_in(w1745), .i_lock(w1747), .o_out(w1746));
	wire w1747;
	repeater #(1, 1'b1, 1, 0) c1747 (.i_clk(tick), .i_in(w199|w297|w517|w737|w957|w1177|w1397|w1617), .i_lock(), .o_out(w1747));
	wire w1952;
	repeater #(1, 1'b1, 0, 0) c1952 (.i_clk(tick), .i_in(w1686|w1696), .i_lock(), .o_out(w1952));
	wire w1959;
	repeater #(1, 1'b1, 0, 0) c1959 (.i_clk(tick), .i_in(w1686|w1696), .i_lock(), .o_out(w1959));
	wire w1964;
	repeater #(1, 1'b1, 1, 0) c1964 (.i_clk(tick), .i_in(w1952), .i_lock(), .o_out(w1964));
	wire w1965;
	repeater #(1, 1'b1, 0, 1) c1965 (.i_clk(tick), .i_in(w1966), .i_lock(w1964), .o_out(w1965));
	wire w1966;
	repeater #(1, 1'b0, 0, 1) c1966 (.i_clk(tick), .i_in(w1965), .i_lock(w1967), .o_out(w1966));
	wire w1967;
	repeater #(1, 1'b1, 1, 0) c1967 (.i_clk(tick), .i_in(w1959), .i_lock(), .o_out(w1967));
	wire w2054;
	repeater #(1, 1'b1, 0, 0) c2054 (.i_clk(tick), .i_in(w1965), .i_lock(), .o_out(w2054));
	wire w2057;
	repeater #(1, 1'b1, 0, 0) c2057 (.i_clk(tick), .i_in(w1965), .i_lock(), .o_out(w2057));
	wire w2184;
	repeater #(1, 1'b1, 1, 0) c2184 (.i_clk(tick), .i_in(w1952|w2054), .i_lock(), .o_out(w2184));
	wire w2185;
	repeater #(1, 1'b1, 0, 1) c2185 (.i_clk(tick), .i_in(w2186), .i_lock(w2184), .o_out(w2185));
	wire w2186;
	repeater #(1, 1'b0, 0, 1) c2186 (.i_clk(tick), .i_in(w2185), .i_lock(w2187), .o_out(w2186));
	wire w2187;
	repeater #(1, 1'b1, 1, 0) c2187 (.i_clk(tick), .i_in(w1959|w2057), .i_lock(), .o_out(w2187));
	wire w2274;
	repeater #(1, 1'b1, 0, 0) c2274 (.i_clk(tick), .i_in(w2185), .i_lock(), .o_out(w2274));
	wire w2277;
	repeater #(1, 1'b1, 0, 0) c2277 (.i_clk(tick), .i_in(w2185), .i_lock(), .o_out(w2277));
	wire w2404;
	repeater #(1, 1'b1, 1, 0) c2404 (.i_clk(tick), .i_in(w1952|w2054|w2274), .i_lock(), .o_out(w2404));
	wire w2405;
	repeater #(1, 1'b1, 0, 1) c2405 (.i_clk(tick), .i_in(w2406), .i_lock(w2404), .o_out(w2405));
	wire w2406;
	repeater #(1, 1'b0, 0, 1) c2406 (.i_clk(tick), .i_in(w2405), .i_lock(w2407), .o_out(w2406));
	wire w2407;
	repeater #(1, 1'b1, 1, 0) c2407 (.i_clk(tick), .i_in(w1959|w2057|w2277), .i_lock(), .o_out(w2407));
	wire w2494;
	repeater #(1, 1'b1, 0, 0) c2494 (.i_clk(tick), .i_in(w2405), .i_lock(), .o_out(w2494));
	wire w2497;
	repeater #(1, 1'b1, 0, 0) c2497 (.i_clk(tick), .i_in(w2405), .i_lock(), .o_out(w2497));
	wire w2624;
	repeater #(1, 1'b1, 1, 0) c2624 (.i_clk(tick), .i_in(w1952|w2054|w2274|w2494), .i_lock(), .o_out(w2624));
	wire w2625;
	repeater #(1, 1'b1, 0, 1) c2625 (.i_clk(tick), .i_in(w2626), .i_lock(w2624), .o_out(w2625));
	wire w2626;
	repeater #(1, 1'b0, 0, 1) c2626 (.i_clk(tick), .i_in(w2625), .i_lock(w2627), .o_out(w2626));
	wire w2627;
	repeater #(1, 1'b1, 1, 0) c2627 (.i_clk(tick), .i_in(w1959|w2057|w2277|w2497), .i_lock(), .o_out(w2627));
	wire w2714;
	repeater #(1, 1'b1, 0, 0) c2714 (.i_clk(tick), .i_in(w2625), .i_lock(), .o_out(w2714));
	wire w2717;
	repeater #(1, 1'b1, 0, 0) c2717 (.i_clk(tick), .i_in(w2625), .i_lock(), .o_out(w2717));
	wire w2844;
	repeater #(1, 1'b1, 1, 0) c2844 (.i_clk(tick), .i_in(w1952|w2054|w2274|w2494|w2714), .i_lock(), .o_out(w2844));
	wire w2845;
	repeater #(1, 1'b1, 0, 1) c2845 (.i_clk(tick), .i_in(w2846), .i_lock(w2844), .o_out(w2845));
	wire w2846;
	repeater #(1, 1'b0, 0, 1) c2846 (.i_clk(tick), .i_in(w2845), .i_lock(w2847), .o_out(w2846));
	wire w2847;
	repeater #(1, 1'b1, 1, 0) c2847 (.i_clk(tick), .i_in(w1959|w2057|w2277|w2497|w2717), .i_lock(), .o_out(w2847));
	wire w2934;
	repeater #(1, 1'b1, 0, 0) c2934 (.i_clk(tick), .i_in(w2845), .i_lock(), .o_out(w2934));
	wire w2937;
	repeater #(1, 1'b1, 0, 0) c2937 (.i_clk(tick), .i_in(w2845), .i_lock(), .o_out(w2937));
	wire w3064;
	repeater #(1, 1'b1, 1, 0) c3064 (.i_clk(tick), .i_in(w1952|w2054|w2274|w2494|w2714|w2934), .i_lock(), .o_out(w3064));
	wire w3065;
	repeater #(1, 1'b1, 0, 1) c3065 (.i_clk(tick), .i_in(w3066), .i_lock(w3064), .o_out(w3065));
	wire w3066;
	repeater #(1, 1'b0, 0, 1) c3066 (.i_clk(tick), .i_in(w3065), .i_lock(w3067), .o_out(w3066));
	wire w3067;
	repeater #(1, 1'b1, 1, 0) c3067 (.i_clk(tick), .i_in(w1959|w2057|w2277|w2497|w2717|w2937), .i_lock(), .o_out(w3067));
	wire w3154;
	repeater #(1, 1'b1, 0, 0) c3154 (.i_clk(tick), .i_in(w3065), .i_lock(), .o_out(w3154));
	wire w3157;
	repeater #(1, 1'b1, 0, 0) c3157 (.i_clk(tick), .i_in(w3065), .i_lock(), .o_out(w3157));
	wire w3284;
	repeater #(1, 1'b1, 1, 0) c3284 (.i_clk(tick), .i_in(w1952|w2054|w2274|w2494|w2714|w2934|w3154), .i_lock(), .o_out(w3284));
	wire w3285;
	repeater #(1, 1'b1, 0, 1) c3285 (.i_clk(tick), .i_in(w3286), .i_lock(w3284), .o_out(w3285));
	wire w3286;
	repeater #(1, 1'b0, 0, 1) c3286 (.i_clk(tick), .i_in(w3285), .i_lock(w3287), .o_out(w3286));
	wire w3287;
	repeater #(1, 1'b1, 1, 0) c3287 (.i_clk(tick), .i_in(w1959|w2057|w2277|w2497|w2717|w2937|w3157), .i_lock(), .o_out(w3287));
	wire w3374;
	repeater #(1, 1'b1, 0, 0) c3374 (.i_clk(tick), .i_in(w3285), .i_lock(), .o_out(w3374));
	wire w3377;
	repeater #(1, 1'b1, 0, 0) c3377 (.i_clk(tick), .i_in(w3285), .i_lock(), .o_out(w3377));
	wire w3445;
	torch #(1'b1) c3445 (.i_clk(tick), .i_in(w3505), .o_out(w3445));
	wire w3446;
	repeater #(2, 1'b0, 0, 0) c3446 (.i_clk(tick), .i_in(w3445), .i_lock(), .o_out(w3446));
	wire w3456;
	repeater #(1, 1'b1, 0, 0) c3456 (.i_clk(tick), .i_in(w3505), .i_lock(), .o_out(w3456));
	wire w3504;
	repeater #(1, 1'b1, 1, 0) c3504 (.i_clk(tick), .i_in(w1952|w2054|w2274|w2494|w2714|w2934|w3154|w3374), .i_lock(), .o_out(w3504));
	wire w3505;
	repeater #(1, 1'b1, 0, 1) c3505 (.i_clk(tick), .i_in(w3506), .i_lock(w3504), .o_out(w3505));
	wire w3506;
	repeater #(1, 1'b0, 0, 1) c3506 (.i_clk(tick), .i_in(w3505), .i_lock(w3507), .o_out(w3506));
	wire w3507;
	repeater #(1, 1'b1, 1, 0) c3507 (.i_clk(tick), .i_in(w1959|w2057|w2277|w2497|w2717|w2937|w3157|w3377), .i_lock(), .o_out(w3507));
	wire w3712;
	repeater #(1, 1'b1, 0, 0) c3712 (.i_clk(tick), .i_in(w3446|w3456), .i_lock(), .o_out(w3712));
	wire w3719;
	repeater #(1, 1'b1, 0, 0) c3719 (.i_clk(tick), .i_in(w3446|w3456), .i_lock(), .o_out(w3719));
	wire w3724;
	repeater #(1, 1'b1, 1, 0) c3724 (.i_clk(tick), .i_in(w3712), .i_lock(), .o_out(w3724));
	wire w3725;
	repeater #(1, 1'b1, 0, 1) c3725 (.i_clk(tick), .i_in(w3726), .i_lock(w3724), .o_out(w3725));
	wire w3726;
	repeater #(1, 1'b0, 0, 1) c3726 (.i_clk(tick), .i_in(w3725), .i_lock(w3727), .o_out(w3726));
	wire w3727;
	repeater #(1, 1'b1, 1, 0) c3727 (.i_clk(tick), .i_in(w3719), .i_lock(), .o_out(w3727));
	wire w3814;
	repeater #(1, 1'b1, 0, 0) c3814 (.i_clk(tick), .i_in(w3725), .i_lock(), .o_out(w3814));
	wire w3817;
	repeater #(1, 1'b1, 0, 0) c3817 (.i_clk(tick), .i_in(w3725), .i_lock(), .o_out(w3817));
	wire w3944;
	repeater #(1, 1'b1, 1, 0) c3944 (.i_clk(tick), .i_in(w3712|w3814), .i_lock(), .o_out(w3944));
	wire w3945;
	repeater #(1, 1'b1, 0, 1) c3945 (.i_clk(tick), .i_in(w3946), .i_lock(w3944), .o_out(w3945));
	wire w3946;
	repeater #(1, 1'b0, 0, 1) c3946 (.i_clk(tick), .i_in(w3945), .i_lock(w3947), .o_out(w3946));
	wire w3947;
	repeater #(1, 1'b1, 1, 0) c3947 (.i_clk(tick), .i_in(w3719|w3817), .i_lock(), .o_out(w3947));
	wire w4034;
	repeater #(1, 1'b1, 0, 0) c4034 (.i_clk(tick), .i_in(w3945), .i_lock(), .o_out(w4034));
	wire w4037;
	repeater #(1, 1'b1, 0, 0) c4037 (.i_clk(tick), .i_in(w3945), .i_lock(), .o_out(w4037));
	wire w4164;
	repeater #(1, 1'b1, 1, 0) c4164 (.i_clk(tick), .i_in(w3712|w3814|w4034), .i_lock(), .o_out(w4164));
	wire w4165;
	repeater #(1, 1'b1, 0, 1) c4165 (.i_clk(tick), .i_in(w4166), .i_lock(w4164), .o_out(w4165));
	wire w4166;
	repeater #(1, 1'b0, 0, 1) c4166 (.i_clk(tick), .i_in(w4165), .i_lock(w4167), .o_out(w4166));
	wire w4167;
	repeater #(1, 1'b1, 1, 0) c4167 (.i_clk(tick), .i_in(w3719|w3817|w4037), .i_lock(), .o_out(w4167));
	wire w4254;
	repeater #(1, 1'b1, 0, 0) c4254 (.i_clk(tick), .i_in(w4165), .i_lock(), .o_out(w4254));
	wire w4257;
	repeater #(1, 1'b1, 0, 0) c4257 (.i_clk(tick), .i_in(w4165), .i_lock(), .o_out(w4257));
	wire w4384;
	repeater #(1, 1'b1, 1, 0) c4384 (.i_clk(tick), .i_in(w3712|w3814|w4034|w4254), .i_lock(), .o_out(w4384));
	wire w4385;
	repeater #(1, 1'b1, 0, 1) c4385 (.i_clk(tick), .i_in(w4386), .i_lock(w4384), .o_out(w4385));
	wire w4386;
	repeater #(1, 1'b0, 0, 1) c4386 (.i_clk(tick), .i_in(w4385), .i_lock(w4387), .o_out(w4386));
	wire w4387;
	repeater #(1, 1'b1, 1, 0) c4387 (.i_clk(tick), .i_in(w3719|w3817|w4037|w4257), .i_lock(), .o_out(w4387));
	wire w4474;
	repeater #(1, 1'b1, 0, 0) c4474 (.i_clk(tick), .i_in(w4385), .i_lock(), .o_out(w4474));
	wire w4477;
	repeater #(1, 1'b1, 0, 0) c4477 (.i_clk(tick), .i_in(w4385), .i_lock(), .o_out(w4477));
	wire w4604;
	repeater #(1, 1'b1, 1, 0) c4604 (.i_clk(tick), .i_in(w3712|w3814|w4034|w4254|w4474), .i_lock(), .o_out(w4604));
	wire w4605;
	repeater #(1, 1'b1, 0, 1) c4605 (.i_clk(tick), .i_in(w4606), .i_lock(w4604), .o_out(w4605));
	wire w4606;
	repeater #(1, 1'b0, 0, 1) c4606 (.i_clk(tick), .i_in(w4605), .i_lock(w4607), .o_out(w4606));
	wire w4607;
	repeater #(1, 1'b1, 1, 0) c4607 (.i_clk(tick), .i_in(w3719|w3817|w4037|w4257|w4477), .i_lock(), .o_out(w4607));
	wire w4694;
	repeater #(1, 1'b1, 0, 0) c4694 (.i_clk(tick), .i_in(w4605), .i_lock(), .o_out(w4694));
	wire w4697;
	repeater #(1, 1'b1, 0, 0) c4697 (.i_clk(tick), .i_in(w4605), .i_lock(), .o_out(w4697));
	wire w4824;
	repeater #(1, 1'b1, 1, 0) c4824 (.i_clk(tick), .i_in(w3712|w3814|w4034|w4254|w4474|w4694), .i_lock(), .o_out(w4824));
	wire w4825;
	repeater #(1, 1'b1, 0, 1) c4825 (.i_clk(tick), .i_in(w4826), .i_lock(w4824), .o_out(w4825));
	wire w4826;
	repeater #(1, 1'b0, 0, 1) c4826 (.i_clk(tick), .i_in(w4825), .i_lock(w4827), .o_out(w4826));
	wire w4827;
	repeater #(1, 1'b1, 1, 0) c4827 (.i_clk(tick), .i_in(w3719|w3817|w4037|w4257|w4477|w4697), .i_lock(), .o_out(w4827));
	wire w4914;
	repeater #(1, 1'b1, 0, 0) c4914 (.i_clk(tick), .i_in(w4825), .i_lock(), .o_out(w4914));
	wire w4917;
	repeater #(1, 1'b1, 0, 0) c4917 (.i_clk(tick), .i_in(w4825), .i_lock(), .o_out(w4917));
	wire w5044;
	repeater #(1, 1'b1, 1, 0) c5044 (.i_clk(tick), .i_in(w3712|w3814|w4034|w4254|w4474|w4694|w4914), .i_lock(), .o_out(w5044));
	wire w5045;
	repeater #(1, 1'b1, 0, 1) c5045 (.i_clk(tick), .i_in(w5046), .i_lock(w5044), .o_out(w5045));
	wire w5046;
	repeater #(1, 1'b0, 0, 1) c5046 (.i_clk(tick), .i_in(w5045), .i_lock(w5047), .o_out(w5046));
	wire w5047;
	repeater #(1, 1'b1, 1, 0) c5047 (.i_clk(tick), .i_in(w3719|w3817|w4037|w4257|w4477|w4697|w4917), .i_lock(), .o_out(w5047));
	wire w5134;
	repeater #(1, 1'b1, 0, 0) c5134 (.i_clk(tick), .i_in(w5045), .i_lock(), .o_out(w5134));
	wire w5137;
	repeater #(1, 1'b0, 0, 0) c5137 (.i_clk(tick), .i_in(w5045), .i_lock(), .o_out(w5137));
	wire w5205;
	torch #(1'b1) c5205 (.i_clk(tick), .i_in(w5265), .o_out(w5205));
	wire w5206;
	repeater #(2, 1'b0, 0, 0) c5206 (.i_clk(tick), .i_in(w5205), .i_lock(), .o_out(w5206));
	wire w5216;
	repeater #(1, 1'b1, 0, 0) c5216 (.i_clk(tick), .i_in(w5265), .i_lock(), .o_out(w5216));
	wire w5264;
	repeater #(1, 1'b1, 1, 0) c5264 (.i_clk(tick), .i_in(w3712|w3814|w4034|w4254|w4474|w4694|w4914|w5134), .i_lock(), .o_out(w5264));
	wire w5265;
	repeater #(1, 1'b1, 0, 1) c5265 (.i_clk(tick), .i_in(w5266), .i_lock(w5264), .o_out(w5265));
	wire w5266;
	repeater #(1, 1'b0, 0, 1) c5266 (.i_clk(tick), .i_in(w5265), .i_lock(w5267), .o_out(w5266));
	wire w5267;
	repeater #(1, 1'b1, 1, 0) c5267 (.i_clk(tick), .i_in(w3719|w3817|w4037|w4257|w4477|w4697|w4917|w5137), .i_lock(), .o_out(w5267));
	wire w5472;
	repeater #(1, 1'b1, 0, 0) c5472 (.i_clk(tick), .i_in(w5206|w5216), .i_lock(), .o_out(w5472));
	wire w5479;
	repeater #(1, 1'b1, 0, 0) c5479 (.i_clk(tick), .i_in(w5206|w5216), .i_lock(), .o_out(w5479));
	wire w5484;
	repeater #(1, 1'b1, 1, 0) c5484 (.i_clk(tick), .i_in(w5472), .i_lock(), .o_out(w5484));
	wire w5485;
	repeater #(1, 1'b1, 0, 1) c5485 (.i_clk(tick), .i_in(w5486), .i_lock(w5484), .o_out(w5485));
	wire w5486;
	repeater #(1, 1'b0, 0, 1) c5486 (.i_clk(tick), .i_in(w5485), .i_lock(w5487), .o_out(w5486));
	wire w5487;
	repeater #(1, 1'b1, 1, 0) c5487 (.i_clk(tick), .i_in(w5479), .i_lock(), .o_out(w5487));
	wire w5566;
	assign outputs[0] = (w5485);
	wire w5574;
	repeater #(1, 1'b1, 0, 0) c5574 (.i_clk(tick), .i_in(w5485), .i_lock(), .o_out(w5574));
	wire w5577;
	repeater #(1, 1'b1, 0, 0) c5577 (.i_clk(tick), .i_in(w5485), .i_lock(), .o_out(w5577));
	wire w5704;
	repeater #(1, 1'b1, 1, 0) c5704 (.i_clk(tick), .i_in(w5472|w5574), .i_lock(), .o_out(w5704));
	wire w5705;
	repeater #(1, 1'b1, 0, 1) c5705 (.i_clk(tick), .i_in(w5706), .i_lock(w5704), .o_out(w5705));
	wire w5706;
	repeater #(1, 1'b0, 0, 1) c5706 (.i_clk(tick), .i_in(w5705), .i_lock(w5707), .o_out(w5706));
	wire w5707;
	repeater #(1, 1'b1, 1, 0) c5707 (.i_clk(tick), .i_in(w5479|w5577), .i_lock(), .o_out(w5707));
	wire w5786;
	assign outputs[1] = (w5705);
	wire w5794;
	repeater #(1, 1'b1, 0, 0) c5794 (.i_clk(tick), .i_in(w5705), .i_lock(), .o_out(w5794));
	wire w5797;
	repeater #(1, 1'b1, 0, 0) c5797 (.i_clk(tick), .i_in(w5705), .i_lock(), .o_out(w5797));
	wire w5924;
	repeater #(1, 1'b1, 1, 0) c5924 (.i_clk(tick), .i_in(w5472|w5574|w5794), .i_lock(), .o_out(w5924));
	wire w5925;
	repeater #(1, 1'b1, 0, 1) c5925 (.i_clk(tick), .i_in(w5926), .i_lock(w5924), .o_out(w5925));
	wire w5926;
	repeater #(1, 1'b0, 0, 1) c5926 (.i_clk(tick), .i_in(w5925), .i_lock(w5927), .o_out(w5926));
	wire w5927;
	repeater #(1, 1'b1, 1, 0) c5927 (.i_clk(tick), .i_in(w5479|w5577|w5797), .i_lock(), .o_out(w5927));
	wire w6006;
	assign outputs[2] = (w5925);
	wire w6014;
	repeater #(1, 1'b1, 0, 0) c6014 (.i_clk(tick), .i_in(w5925), .i_lock(), .o_out(w6014));
	wire w6017;
	repeater #(1, 1'b1, 0, 0) c6017 (.i_clk(tick), .i_in(w5925), .i_lock(), .o_out(w6017));
	wire w6144;
	repeater #(1, 1'b1, 1, 0) c6144 (.i_clk(tick), .i_in(w5472|w5574|w5794|w6014), .i_lock(), .o_out(w6144));
	wire w6145;
	repeater #(1, 1'b1, 0, 1) c6145 (.i_clk(tick), .i_in(w6146), .i_lock(w6144), .o_out(w6145));
	wire w6146;
	repeater #(1, 1'b0, 0, 1) c6146 (.i_clk(tick), .i_in(w6145), .i_lock(w6147), .o_out(w6146));
	wire w6147;
	repeater #(1, 1'b1, 1, 0) c6147 (.i_clk(tick), .i_in(w5479|w5577|w5797|w6017), .i_lock(), .o_out(w6147));
	wire w6226;
	assign outputs[3] = (w6145);
	wire w6234;
	repeater #(1, 1'b1, 0, 0) c6234 (.i_clk(tick), .i_in(w6145), .i_lock(), .o_out(w6234));
	wire w6237;
	repeater #(1, 1'b1, 0, 0) c6237 (.i_clk(tick), .i_in(w6145), .i_lock(), .o_out(w6237));
	wire w6364;
	repeater #(1, 1'b1, 1, 0) c6364 (.i_clk(tick), .i_in(w5472|w5574|w5794|w6014|w6234), .i_lock(), .o_out(w6364));
	wire w6365;
	repeater #(1, 1'b1, 0, 1) c6365 (.i_clk(tick), .i_in(w6366), .i_lock(w6364), .o_out(w6365));
	wire w6366;
	repeater #(1, 1'b0, 0, 1) c6366 (.i_clk(tick), .i_in(w6365), .i_lock(w6367), .o_out(w6366));
	wire w6367;
	repeater #(1, 1'b1, 1, 0) c6367 (.i_clk(tick), .i_in(w5479|w5577|w5797|w6017|w6237), .i_lock(), .o_out(w6367));
	wire w6446;
	assign outputs[4] = (w6365);
	wire w6454;
	repeater #(1, 1'b1, 0, 0) c6454 (.i_clk(tick), .i_in(w6365), .i_lock(), .o_out(w6454));
	wire w6457;
	repeater #(1, 1'b1, 0, 0) c6457 (.i_clk(tick), .i_in(w6365), .i_lock(), .o_out(w6457));
	wire w6584;
	repeater #(1, 1'b1, 1, 0) c6584 (.i_clk(tick), .i_in(w5472|w5574|w5794|w6014|w6234|w6454), .i_lock(), .o_out(w6584));
	wire w6585;
	repeater #(1, 1'b1, 0, 1) c6585 (.i_clk(tick), .i_in(w6586), .i_lock(w6584), .o_out(w6585));
	wire w6586;
	repeater #(1, 1'b0, 0, 1) c6586 (.i_clk(tick), .i_in(w6585), .i_lock(w6587), .o_out(w6586));
	wire w6587;
	repeater #(1, 1'b1, 1, 0) c6587 (.i_clk(tick), .i_in(w5479|w5577|w5797|w6017|w6237|w6457), .i_lock(), .o_out(w6587));
	wire w6666;
	assign outputs[5] = (w6585);
	wire w6674;
	repeater #(1, 1'b1, 0, 0) c6674 (.i_clk(tick), .i_in(w6585), .i_lock(), .o_out(w6674));
	wire w6677;
	repeater #(1, 1'b1, 0, 0) c6677 (.i_clk(tick), .i_in(w6585), .i_lock(), .o_out(w6677));
	wire w6804;
	repeater #(1, 1'b1, 1, 0) c6804 (.i_clk(tick), .i_in(w5472|w5574|w5794|w6014|w6234|w6454|w6674), .i_lock(), .o_out(w6804));
	wire w6805;
	repeater #(1, 1'b1, 0, 1) c6805 (.i_clk(tick), .i_in(w6806), .i_lock(w6804), .o_out(w6805));
	wire w6806;
	repeater #(1, 1'b0, 0, 1) c6806 (.i_clk(tick), .i_in(w6805), .i_lock(w6807), .o_out(w6806));
	wire w6807;
	repeater #(1, 1'b1, 1, 0) c6807 (.i_clk(tick), .i_in(w5479|w5577|w5797|w6017|w6237|w6457|w6677), .i_lock(), .o_out(w6807));
	wire w6886;
	assign outputs[6] = (w6805);
	wire w6894;
	repeater #(1, 1'b1, 0, 0) c6894 (.i_clk(tick), .i_in(w6805), .i_lock(), .o_out(w6894));
	wire w6897;
	repeater #(1, 1'b1, 0, 0) c6897 (.i_clk(tick), .i_in(w6805), .i_lock(), .o_out(w6897));
	wire w7024;
	repeater #(1, 1'b1, 1, 0) c7024 (.i_clk(tick), .i_in(w5472|w5574|w5794|w6014|w6234|w6454|w6674|w6894), .i_lock(), .o_out(w7024));
	wire w7025;
	repeater #(1, 1'b1, 0, 1) c7025 (.i_clk(tick), .i_in(w7026), .i_lock(w7024), .o_out(w7025));
	wire w7026;
	repeater #(1, 1'b0, 0, 1) c7026 (.i_clk(tick), .i_in(w7025), .i_lock(w7027), .o_out(w7026));
	wire w7027;
	repeater #(1, 1'b1, 1, 0) c7027 (.i_clk(tick), .i_in(w5479|w5577|w5797|w6017|w6237|w6457|w6677|w6897), .i_lock(), .o_out(w7027));
	wire w7106;
	assign outputs[7] = (w7025);
endmodule