parameter num_outputs = 32;
parameter num_inputs = 1;
parameter num_bytes = 8'd4;