// EBAB.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module EBAB (
		input  wire        clk_clk,                    //                  clk.clk
		input  wire [11:0] ebab_address,               //                 ebab.address
		input  wire [1:0]  ebab_byte_enable,           //                     .byte_enable
		input  wire        ebab_read,                  //                     .read
		input  wire        ebab_write,                 //                     .write
		input  wire [15:0] ebab_write_data,            //                     .write_data
		output wire        ebab_acknowledge,           //                     .acknowledge
		output wire [15:0] ebab_read_data,             //                     .read_data
		output wire        hps_io_reset_n,             //               hps_io.reset_n
		input  wire        reset_reset_n,              //                reset.reset_n
		output wire        sdram_clk_clk,              //            sdram_clk.clk
		input  wire        system_pll_ref_clk_clk,     //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset  // system_pll_ref_reset.reset
	);

	wire         pll_sys_clk_clk;                // PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, EBAB:clk, rst_controller:clk]
	wire  [31:0] arm_a9_hps_f2h_irq0_irq;        // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;        // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         rst_controller_reset_out_reset; // rst_controller:reset_out -> EBAB:reset
	wire         pll_reset_source_reset;         // PLL:reset_source_reset -> rst_controller:reset_in0

	EBAB_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a          (),                        //            memory.mem_a
		.mem_ba         (),                        //                  .mem_ba
		.mem_ck         (),                        //                  .mem_ck
		.mem_ck_n       (),                        //                  .mem_ck_n
		.mem_cke        (),                        //                  .mem_cke
		.mem_cs_n       (),                        //                  .mem_cs_n
		.mem_ras_n      (),                        //                  .mem_ras_n
		.mem_cas_n      (),                        //                  .mem_cas_n
		.mem_we_n       (),                        //                  .mem_we_n
		.mem_reset_n    (),                        //                  .mem_reset_n
		.mem_dq         (),                        //                  .mem_dq
		.mem_dqs        (),                        //                  .mem_dqs
		.mem_dqs_n      (),                        //                  .mem_dqs_n
		.mem_odt        (),                        //                  .mem_odt
		.mem_dm         (),                        //                  .mem_dm
		.oct_rzqin      (),                        //                  .oct_rzqin
		.h2f_rst_n      (hps_io_reset_n),          //         h2f_reset.reset_n
		.h2f_axi_clk    (pll_sys_clk_clk),         //     h2f_axi_clock.clk
		.h2f_AWID       (),                        //    h2f_axi_master.awid
		.h2f_AWADDR     (),                        //                  .awaddr
		.h2f_AWLEN      (),                        //                  .awlen
		.h2f_AWSIZE     (),                        //                  .awsize
		.h2f_AWBURST    (),                        //                  .awburst
		.h2f_AWLOCK     (),                        //                  .awlock
		.h2f_AWCACHE    (),                        //                  .awcache
		.h2f_AWPROT     (),                        //                  .awprot
		.h2f_AWVALID    (),                        //                  .awvalid
		.h2f_AWREADY    (),                        //                  .awready
		.h2f_WID        (),                        //                  .wid
		.h2f_WDATA      (),                        //                  .wdata
		.h2f_WSTRB      (),                        //                  .wstrb
		.h2f_WLAST      (),                        //                  .wlast
		.h2f_WVALID     (),                        //                  .wvalid
		.h2f_WREADY     (),                        //                  .wready
		.h2f_BID        (),                        //                  .bid
		.h2f_BRESP      (),                        //                  .bresp
		.h2f_BVALID     (),                        //                  .bvalid
		.h2f_BREADY     (),                        //                  .bready
		.h2f_ARID       (),                        //                  .arid
		.h2f_ARADDR     (),                        //                  .araddr
		.h2f_ARLEN      (),                        //                  .arlen
		.h2f_ARSIZE     (),                        //                  .arsize
		.h2f_ARBURST    (),                        //                  .arburst
		.h2f_ARLOCK     (),                        //                  .arlock
		.h2f_ARCACHE    (),                        //                  .arcache
		.h2f_ARPROT     (),                        //                  .arprot
		.h2f_ARVALID    (),                        //                  .arvalid
		.h2f_ARREADY    (),                        //                  .arready
		.h2f_RID        (),                        //                  .rid
		.h2f_RDATA      (),                        //                  .rdata
		.h2f_RRESP      (),                        //                  .rresp
		.h2f_RLAST      (),                        //                  .rlast
		.h2f_RVALID     (),                        //                  .rvalid
		.h2f_RREADY     (),                        //                  .rready
		.f2h_axi_clk    (pll_sys_clk_clk),         //     f2h_axi_clock.clk
		.f2h_AWID       (),                        //     f2h_axi_slave.awid
		.f2h_AWADDR     (),                        //                  .awaddr
		.f2h_AWLEN      (),                        //                  .awlen
		.f2h_AWSIZE     (),                        //                  .awsize
		.f2h_AWBURST    (),                        //                  .awburst
		.f2h_AWLOCK     (),                        //                  .awlock
		.f2h_AWCACHE    (),                        //                  .awcache
		.f2h_AWPROT     (),                        //                  .awprot
		.f2h_AWVALID    (),                        //                  .awvalid
		.f2h_AWREADY    (),                        //                  .awready
		.f2h_AWUSER     (),                        //                  .awuser
		.f2h_WID        (),                        //                  .wid
		.f2h_WDATA      (),                        //                  .wdata
		.f2h_WSTRB      (),                        //                  .wstrb
		.f2h_WLAST      (),                        //                  .wlast
		.f2h_WVALID     (),                        //                  .wvalid
		.f2h_WREADY     (),                        //                  .wready
		.f2h_BID        (),                        //                  .bid
		.f2h_BRESP      (),                        //                  .bresp
		.f2h_BVALID     (),                        //                  .bvalid
		.f2h_BREADY     (),                        //                  .bready
		.f2h_ARID       (),                        //                  .arid
		.f2h_ARADDR     (),                        //                  .araddr
		.f2h_ARLEN      (),                        //                  .arlen
		.f2h_ARSIZE     (),                        //                  .arsize
		.f2h_ARBURST    (),                        //                  .arburst
		.f2h_ARLOCK     (),                        //                  .arlock
		.f2h_ARCACHE    (),                        //                  .arcache
		.f2h_ARPROT     (),                        //                  .arprot
		.f2h_ARVALID    (),                        //                  .arvalid
		.f2h_ARREADY    (),                        //                  .arready
		.f2h_ARUSER     (),                        //                  .aruser
		.f2h_RID        (),                        //                  .rid
		.f2h_RDATA      (),                        //                  .rdata
		.f2h_RRESP      (),                        //                  .rresp
		.f2h_RLAST      (),                        //                  .rlast
		.f2h_RVALID     (),                        //                  .rvalid
		.f2h_RREADY     (),                        //                  .rready
		.h2f_lw_axi_clk (pll_sys_clk_clk),         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (),                        // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (),                        //                  .awaddr
		.h2f_lw_AWLEN   (),                        //                  .awlen
		.h2f_lw_AWSIZE  (),                        //                  .awsize
		.h2f_lw_AWBURST (),                        //                  .awburst
		.h2f_lw_AWLOCK  (),                        //                  .awlock
		.h2f_lw_AWCACHE (),                        //                  .awcache
		.h2f_lw_AWPROT  (),                        //                  .awprot
		.h2f_lw_AWVALID (),                        //                  .awvalid
		.h2f_lw_AWREADY (),                        //                  .awready
		.h2f_lw_WID     (),                        //                  .wid
		.h2f_lw_WDATA   (),                        //                  .wdata
		.h2f_lw_WSTRB   (),                        //                  .wstrb
		.h2f_lw_WLAST   (),                        //                  .wlast
		.h2f_lw_WVALID  (),                        //                  .wvalid
		.h2f_lw_WREADY  (),                        //                  .wready
		.h2f_lw_BID     (),                        //                  .bid
		.h2f_lw_BRESP   (),                        //                  .bresp
		.h2f_lw_BVALID  (),                        //                  .bvalid
		.h2f_lw_BREADY  (),                        //                  .bready
		.h2f_lw_ARID    (),                        //                  .arid
		.h2f_lw_ARADDR  (),                        //                  .araddr
		.h2f_lw_ARLEN   (),                        //                  .arlen
		.h2f_lw_ARSIZE  (),                        //                  .arsize
		.h2f_lw_ARBURST (),                        //                  .arburst
		.h2f_lw_ARLOCK  (),                        //                  .arlock
		.h2f_lw_ARCACHE (),                        //                  .arcache
		.h2f_lw_ARPROT  (),                        //                  .arprot
		.h2f_lw_ARVALID (),                        //                  .arvalid
		.h2f_lw_ARREADY (),                        //                  .arready
		.h2f_lw_RID     (),                        //                  .rid
		.h2f_lw_RDATA   (),                        //                  .rdata
		.h2f_lw_RRESP   (),                        //                  .rresp
		.h2f_lw_RLAST   (),                        //                  .rlast
		.h2f_lw_RVALID  (),                        //                  .rvalid
		.h2f_lw_RREADY  (),                        //                  .rready
		.f2h_irq_p0     (arm_a9_hps_f2h_irq0_irq), //          f2h_irq0.irq
		.f2h_irq_p1     (arm_a9_hps_f2h_irq1_irq)  //          f2h_irq1.irq
	);

	EBAB_EBAB ebab (
		.clk                (pll_sys_clk_clk),                //                clk.clk
		.reset              (rst_controller_reset_out_reset), //              reset.reset
		.avalon_readdata    (),                               //      avalon_master.readdata
		.avalon_waitrequest (),                               //                   .waitrequest
		.avalon_byteenable  (),                               //                   .byteenable
		.avalon_read        (),                               //                   .read
		.avalon_write       (),                               //                   .write
		.avalon_writedata   (),                               //                   .writedata
		.avalon_address     (),                               //                   .address
		.address            (ebab_address),                   // external_interface.export
		.byte_enable        (ebab_byte_enable),               //                   .export
		.read               (ebab_read),                      //                   .export
		.write              (ebab_write),                     //                   .export
		.write_data         (ebab_write_data),                //                   .export
		.acknowledge        (ebab_acknowledge),               //                   .export
		.read_data          (ebab_read_data)                  //                   .export
	);

	EBAB_PLL pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),     //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset), //    ref_reset.reset
		.sys_clk_clk        (pll_sys_clk_clk),            //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),              //    sdram_clk.clk
		.reset_source_reset (pll_reset_source_reset)      // reset_source.reset
	);

	EBAB_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq0_irq)  //    sender.irq
	);

	EBAB_irq_mapper irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (pll_reset_source_reset),         // reset_in0.reset
		.clk            (pll_sys_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
